-- eth_std_main_system_ethernet_subsystem.vhd

-- Generated using ACDS version 16.1 196

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity eth_std_main_system_ethernet_subsystem is
	port (
		descriptor_memory_s2_address     : in  std_logic_vector(10 downto 0) := (others => '0'); --     descriptor_memory_s2.address
		descriptor_memory_s2_chipselect  : in  std_logic                     := '0';             --                         .chipselect
		descriptor_memory_s2_clken       : in  std_logic                     := '0';             --                         .clken
		descriptor_memory_s2_write       : in  std_logic                     := '0';             --                         .write
		descriptor_memory_s2_readdata    : out std_logic_vector(31 downto 0);                    --                         .readdata
		descriptor_memory_s2_writedata   : in  std_logic_vector(31 downto 0) := (others => '0'); --                         .writedata
		descriptor_memory_s2_byteenable  : in  std_logic_vector(3 downto 0)  := (others => '0'); --                         .byteenable
		ethernet_bridge_s0_waitrequest   : out std_logic;                                        --       ethernet_bridge_s0.waitrequest
		ethernet_bridge_s0_readdata      : out std_logic_vector(31 downto 0);                    --                         .readdata
		ethernet_bridge_s0_readdatavalid : out std_logic;                                        --                         .readdatavalid
		ethernet_bridge_s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => '0'); --                         .burstcount
		ethernet_bridge_s0_writedata     : in  std_logic_vector(31 downto 0) := (others => '0'); --                         .writedata
		ethernet_bridge_s0_address       : in  std_logic_vector(10 downto 0) := (others => '0'); --                         .address
		ethernet_bridge_s0_write         : in  std_logic                     := '0';             --                         .write
		ethernet_bridge_s0_read          : in  std_logic                     := '0';             --                         .read
		ethernet_bridge_s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => '0'); --                         .byteenable
		ethernet_bridge_s0_debugaccess   : in  std_logic                     := '0';             --                         .debugaccess
		ethernet_subsys_clk_in_clk       : in  std_logic                     := '0';             --   ethernet_subsys_clk_in.clk
		ethernet_subsys_reset_in_reset_n : in  std_logic                     := '0';             -- ethernet_subsys_reset_in.reset_n
		mac_gmii_connection_gmii_rx_d    : in  std_logic_vector(7 downto 0)  := (others => '0'); --      mac_gmii_connection.gmii_rx_d
		mac_gmii_connection_gmii_rx_dv   : in  std_logic                     := '0';             --                         .gmii_rx_dv
		mac_gmii_connection_gmii_rx_err  : in  std_logic                     := '0';             --                         .gmii_rx_err
		mac_gmii_connection_gmii_tx_d    : out std_logic_vector(7 downto 0);                     --                         .gmii_tx_d
		mac_gmii_connection_gmii_tx_en   : out std_logic;                                        --                         .gmii_tx_en
		mac_gmii_connection_gmii_tx_err  : out std_logic;                                        --                         .gmii_tx_err
		mac_mdio_connection_mdc          : out std_logic;                                        --      mac_mdio_connection.mdc
		mac_mdio_connection_mdio_in      : in  std_logic                     := '0';             --                         .mdio_in
		mac_mdio_connection_mdio_out     : out std_logic;                                        --                         .mdio_out
		mac_mdio_connection_mdio_oen     : out std_logic;                                        --                         .mdio_oen
		mac_mii_connection_mii_rx_d      : in  std_logic_vector(3 downto 0)  := (others => '0'); --       mac_mii_connection.mii_rx_d
		mac_mii_connection_mii_rx_dv     : in  std_logic                     := '0';             --                         .mii_rx_dv
		mac_mii_connection_mii_rx_err    : in  std_logic                     := '0';             --                         .mii_rx_err
		mac_mii_connection_mii_tx_d      : out std_logic_vector(3 downto 0);                     --                         .mii_tx_d
		mac_mii_connection_mii_tx_en     : out std_logic;                                        --                         .mii_tx_en
		mac_mii_connection_mii_tx_err    : out std_logic;                                        --                         .mii_tx_err
		mac_mii_connection_mii_crs       : in  std_logic                     := '0';             --                         .mii_crs
		mac_mii_connection_mii_col       : in  std_logic                     := '0';             --                         .mii_col
		mac_status_connection_set_10     : in  std_logic                     := '0';             --    mac_status_connection.set_10
		mac_status_connection_set_1000   : in  std_logic                     := '0';             --                         .set_1000
		mac_status_connection_eth_mode   : out std_logic;                                        --                         .eth_mode
		mac_status_connection_ena_10     : out std_logic;                                        --                         .ena_10
		misc_connection_xon_gen          : in  std_logic                     := '0';             --          misc_connection.xon_gen
		misc_connection_xoff_gen         : in  std_logic                     := '0';             --                         .xoff_gen
		misc_connection_ff_tx_crc_fwd    : in  std_logic                     := '0';             --                         .ff_tx_crc_fwd
		misc_connection_ff_tx_septy      : out std_logic;                                        --                         .ff_tx_septy
		misc_connection_tx_ff_uflow      : out std_logic;                                        --                         .tx_ff_uflow
		misc_connection_ff_tx_a_full     : out std_logic;                                        --                         .ff_tx_a_full
		misc_connection_ff_tx_a_empty    : out std_logic;                                        --                         .ff_tx_a_empty
		misc_connection_rx_err_stat      : out std_logic_vector(17 downto 0);                    --                         .rx_err_stat
		misc_connection_rx_frm_type      : out std_logic_vector(3 downto 0);                     --                         .rx_frm_type
		misc_connection_ff_rx_dsav       : out std_logic;                                        --                         .ff_rx_dsav
		misc_connection_ff_rx_a_full     : out std_logic;                                        --                         .ff_rx_a_full
		misc_connection_ff_rx_a_empty    : out std_logic;                                        --                         .ff_rx_a_empty
		rx_clock_clk                     : in  std_logic                     := '0';             --                 rx_clock.clk
		sgdma_bridge_m0_waitrequest      : in  std_logic                     := '0';             --          sgdma_bridge_m0.waitrequest
		sgdma_bridge_m0_readdata         : in  std_logic_vector(31 downto 0) := (others => '0'); --                         .readdata
		sgdma_bridge_m0_readdatavalid    : in  std_logic                     := '0';             --                         .readdatavalid
		sgdma_bridge_m0_burstcount       : out std_logic_vector(0 downto 0);                     --                         .burstcount
		sgdma_bridge_m0_writedata        : out std_logic_vector(31 downto 0);                    --                         .writedata
		sgdma_bridge_m0_address          : out std_logic_vector(30 downto 0);                    --                         .address
		sgdma_bridge_m0_write            : out std_logic;                                        --                         .write
		sgdma_bridge_m0_read             : out std_logic;                                        --                         .read
		sgdma_bridge_m0_byteenable       : out std_logic_vector(3 downto 0);                     --                         .byteenable
		sgdma_bridge_m0_debugaccess      : out std_logic;                                        --                         .debugaccess
		sgdma_rx_csr_irq_irq             : out std_logic;                                        --         sgdma_rx_csr_irq.irq
		sgdma_tx_csr_irq_irq             : out std_logic;                                        --         sgdma_tx_csr_irq.irq
		tx_clock_clk                     : in  std_logic                     := '0'              --                 tx_clock.clk
	);
end entity eth_std_main_system_ethernet_subsystem;

architecture rtl of eth_std_main_system_ethernet_subsystem is
	component eth_std_main_system_ethernet_subsystem_descriptor_memory is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			address     : in  std_logic_vector(10 downto 0) := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			address2    : in  std_logic_vector(10 downto 0) := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk2        : in  std_logic                     := 'X';             -- clk
			reset2      : in  std_logic                     := 'X';             -- reset
			reset_req2  : in  std_logic                     := 'X';             -- reset_req
			freeze      : in  std_logic                     := 'X'              -- freeze
		);
	end component eth_std_main_system_ethernet_subsystem_descriptor_memory;

	component eth_std_main_system_ethernet_subsystem_sgdma_rx is
		port (
			clk                           : in  std_logic                     := 'X';             -- clk
			system_reset_n                : in  std_logic                     := 'X';             -- reset_n
			csr_chipselect                : in  std_logic                     := 'X';             -- chipselect
			csr_address                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			csr_read                      : in  std_logic                     := 'X';             -- read
			csr_write                     : in  std_logic                     := 'X';             -- write
			csr_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			csr_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			descriptor_read_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			descriptor_read_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			descriptor_read_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			descriptor_read_address       : out std_logic_vector(31 downto 0);                    -- address
			descriptor_read_read          : out std_logic;                                        -- read
			descriptor_write_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			descriptor_write_address      : out std_logic_vector(31 downto 0);                    -- address
			descriptor_write_write        : out std_logic;                                        -- write
			descriptor_write_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			csr_irq                       : out std_logic;                                        -- irq
			in_startofpacket              : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket                : in  std_logic                     := 'X';             -- endofpacket
			in_data                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_valid                      : in  std_logic                     := 'X';             -- valid
			in_ready                      : out std_logic;                                        -- ready
			in_empty                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			in_error                      : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- error
			m_write_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			m_write_address               : out std_logic_vector(31 downto 0);                    -- address
			m_write_write                 : out std_logic;                                        -- write
			m_write_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			m_write_byteenable            : out std_logic_vector(3 downto 0)                      -- byteenable
		);
	end component eth_std_main_system_ethernet_subsystem_sgdma_rx;

	component eth_std_main_system_ethernet_subsystem_sgdma_tx is
		port (
			clk                           : in  std_logic                     := 'X';             -- clk
			system_reset_n                : in  std_logic                     := 'X';             -- reset_n
			csr_chipselect                : in  std_logic                     := 'X';             -- chipselect
			csr_address                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			csr_read                      : in  std_logic                     := 'X';             -- read
			csr_write                     : in  std_logic                     := 'X';             -- write
			csr_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			csr_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			descriptor_read_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			descriptor_read_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			descriptor_read_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			descriptor_read_address       : out std_logic_vector(31 downto 0);                    -- address
			descriptor_read_read          : out std_logic;                                        -- read
			descriptor_write_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			descriptor_write_address      : out std_logic_vector(31 downto 0);                    -- address
			descriptor_write_write        : out std_logic;                                        -- write
			descriptor_write_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			csr_irq                       : out std_logic;                                        -- irq
			m_read_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m_read_readdatavalid          : in  std_logic                     := 'X';             -- readdatavalid
			m_read_waitrequest            : in  std_logic                     := 'X';             -- waitrequest
			m_read_address                : out std_logic_vector(31 downto 0);                    -- address
			m_read_read                   : out std_logic;                                        -- read
			out_data                      : out std_logic_vector(31 downto 0);                    -- data
			out_valid                     : out std_logic;                                        -- valid
			out_ready                     : in  std_logic                     := 'X';             -- ready
			out_endofpacket               : out std_logic;                                        -- endofpacket
			out_startofpacket             : out std_logic;                                        -- startofpacket
			out_empty                     : out std_logic_vector(1 downto 0);                     -- empty
			out_error                     : out std_logic                                         -- error
		);
	end component eth_std_main_system_ethernet_subsystem_sgdma_tx;

	component eth_std_main_system_ethernet_subsystem_tse_mac is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			reg_addr      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			reg_data_out  : out std_logic_vector(31 downto 0);                    -- readdata
			reg_rd        : in  std_logic                     := 'X';             -- read
			reg_data_in   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			reg_wr        : in  std_logic                     := 'X';             -- write
			reg_busy      : out std_logic;                                        -- waitrequest
			tx_clk        : in  std_logic                     := 'X';             -- clk
			rx_clk        : in  std_logic                     := 'X';             -- clk
			set_10        : in  std_logic                     := 'X';             -- set_10
			set_1000      : in  std_logic                     := 'X';             -- set_1000
			eth_mode      : out std_logic;                                        -- eth_mode
			ena_10        : out std_logic;                                        -- ena_10
			gm_rx_d       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- gmii_rx_d
			gm_rx_dv      : in  std_logic                     := 'X';             -- gmii_rx_dv
			gm_rx_err     : in  std_logic                     := 'X';             -- gmii_rx_err
			gm_tx_d       : out std_logic_vector(7 downto 0);                     -- gmii_tx_d
			gm_tx_en      : out std_logic;                                        -- gmii_tx_en
			gm_tx_err     : out std_logic;                                        -- gmii_tx_err
			m_rx_d        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- mii_rx_d
			m_rx_en       : in  std_logic                     := 'X';             -- mii_rx_dv
			m_rx_err      : in  std_logic                     := 'X';             -- mii_rx_err
			m_tx_d        : out std_logic_vector(3 downto 0);                     -- mii_tx_d
			m_tx_en       : out std_logic;                                        -- mii_tx_en
			m_tx_err      : out std_logic;                                        -- mii_tx_err
			m_rx_crs      : in  std_logic                     := 'X';             -- mii_crs
			m_rx_col      : in  std_logic                     := 'X';             -- mii_col
			ff_rx_clk     : in  std_logic                     := 'X';             -- clk
			ff_tx_clk     : in  std_logic                     := 'X';             -- clk
			ff_rx_data    : out std_logic_vector(31 downto 0);                    -- data
			ff_rx_eop     : out std_logic;                                        -- endofpacket
			rx_err        : out std_logic_vector(5 downto 0);                     -- error
			ff_rx_mod     : out std_logic_vector(1 downto 0);                     -- empty
			ff_rx_rdy     : in  std_logic                     := 'X';             -- ready
			ff_rx_sop     : out std_logic;                                        -- startofpacket
			ff_rx_dval    : out std_logic;                                        -- valid
			ff_tx_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			ff_tx_eop     : in  std_logic                     := 'X';             -- endofpacket
			ff_tx_err     : in  std_logic                     := 'X';             -- error
			ff_tx_mod     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			ff_tx_rdy     : out std_logic;                                        -- ready
			ff_tx_sop     : in  std_logic                     := 'X';             -- startofpacket
			ff_tx_wren    : in  std_logic                     := 'X';             -- valid
			mdc           : out std_logic;                                        -- mdc
			mdio_in       : in  std_logic                     := 'X';             -- mdio_in
			mdio_out      : out std_logic;                                        -- mdio_out
			mdio_oen      : out std_logic;                                        -- mdio_oen
			xon_gen       : in  std_logic                     := 'X';             -- xon_gen
			xoff_gen      : in  std_logic                     := 'X';             -- xoff_gen
			ff_tx_crc_fwd : in  std_logic                     := 'X';             -- ff_tx_crc_fwd
			ff_tx_septy   : out std_logic;                                        -- ff_tx_septy
			tx_ff_uflow   : out std_logic;                                        -- tx_ff_uflow
			ff_tx_a_full  : out std_logic;                                        -- ff_tx_a_full
			ff_tx_a_empty : out std_logic;                                        -- ff_tx_a_empty
			rx_err_stat   : out std_logic_vector(17 downto 0);                    -- rx_err_stat
			rx_frm_type   : out std_logic_vector(3 downto 0);                     -- rx_frm_type
			ff_rx_dsav    : out std_logic;                                        -- ff_rx_dsav
			ff_rx_a_full  : out std_logic;                                        -- ff_rx_a_full
			ff_rx_a_empty : out std_logic                                         -- ff_rx_a_empty
		);
	end component eth_std_main_system_ethernet_subsystem_tse_mac;

	component eth_std_main_system_ethernet_subsystem_mm_interconnect_0 is
		port (
			clk_clk_clk                                : in  std_logic                     := 'X';             -- clk
			sgdma_tx_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			sgdma_rx_descriptor_read_address           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_rx_descriptor_read_waitrequest       : out std_logic;                                        -- waitrequest
			sgdma_rx_descriptor_read_read              : in  std_logic                     := 'X';             -- read
			sgdma_rx_descriptor_read_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			sgdma_rx_descriptor_read_readdatavalid     : out std_logic;                                        -- readdatavalid
			sgdma_rx_descriptor_write_address          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_rx_descriptor_write_waitrequest      : out std_logic;                                        -- waitrequest
			sgdma_rx_descriptor_write_write            : in  std_logic                     := 'X';             -- write
			sgdma_rx_descriptor_write_writedata        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			sgdma_tx_descriptor_read_address           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_tx_descriptor_read_waitrequest       : out std_logic;                                        -- waitrequest
			sgdma_tx_descriptor_read_read              : in  std_logic                     := 'X';             -- read
			sgdma_tx_descriptor_read_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			sgdma_tx_descriptor_read_readdatavalid     : out std_logic;                                        -- readdatavalid
			sgdma_tx_descriptor_write_address          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_tx_descriptor_write_waitrequest      : out std_logic;                                        -- waitrequest
			sgdma_tx_descriptor_write_write            : in  std_logic                     := 'X';             -- write
			sgdma_tx_descriptor_write_writedata        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			descriptor_memory_s1_address               : out std_logic_vector(10 downto 0);                    -- address
			descriptor_memory_s1_write                 : out std_logic;                                        -- write
			descriptor_memory_s1_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			descriptor_memory_s1_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			descriptor_memory_s1_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			descriptor_memory_s1_chipselect            : out std_logic;                                        -- chipselect
			descriptor_memory_s1_clken                 : out std_logic                                         -- clken
		);
	end component eth_std_main_system_ethernet_subsystem_mm_interconnect_0;

	component eth_std_main_system_ethernet_subsystem_mm_interconnect_1 is
		port (
			clk_clk_clk                                       : in  std_logic                     := 'X';             -- clk
			ethernet_bridge_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			ethernet_bridge_m0_address                        : in  std_logic_vector(10 downto 0) := (others => 'X'); -- address
			ethernet_bridge_m0_waitrequest                    : out std_logic;                                        -- waitrequest
			ethernet_bridge_m0_burstcount                     : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			ethernet_bridge_m0_byteenable                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			ethernet_bridge_m0_read                           : in  std_logic                     := 'X';             -- read
			ethernet_bridge_m0_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			ethernet_bridge_m0_readdatavalid                  : out std_logic;                                        -- readdatavalid
			ethernet_bridge_m0_write                          : in  std_logic                     := 'X';             -- write
			ethernet_bridge_m0_writedata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			ethernet_bridge_m0_debugaccess                    : in  std_logic                     := 'X';             -- debugaccess
			sgdma_rx_csr_address                              : out std_logic_vector(3 downto 0);                     -- address
			sgdma_rx_csr_write                                : out std_logic;                                        -- write
			sgdma_rx_csr_read                                 : out std_logic;                                        -- read
			sgdma_rx_csr_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sgdma_rx_csr_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			sgdma_rx_csr_chipselect                           : out std_logic;                                        -- chipselect
			sgdma_tx_csr_address                              : out std_logic_vector(3 downto 0);                     -- address
			sgdma_tx_csr_write                                : out std_logic;                                        -- write
			sgdma_tx_csr_read                                 : out std_logic;                                        -- read
			sgdma_tx_csr_readdata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sgdma_tx_csr_writedata                            : out std_logic_vector(31 downto 0);                    -- writedata
			sgdma_tx_csr_chipselect                           : out std_logic;                                        -- chipselect
			tse_mac_control_port_address                      : out std_logic_vector(7 downto 0);                     -- address
			tse_mac_control_port_write                        : out std_logic;                                        -- write
			tse_mac_control_port_read                         : out std_logic;                                        -- read
			tse_mac_control_port_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			tse_mac_control_port_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			tse_mac_control_port_waitrequest                  : in  std_logic                     := 'X'              -- waitrequest
		);
	end component eth_std_main_system_ethernet_subsystem_mm_interconnect_1;

	component eth_std_main_system_ethernet_subsystem_mm_interconnect_2 is
		port (
			clk_clk_clk                                : in  std_logic                     := 'X';             -- clk
			sgdma_tx_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			sgdma_rx_m_write_address                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_rx_m_write_waitrequest               : out std_logic;                                        -- waitrequest
			sgdma_rx_m_write_byteenable                : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			sgdma_rx_m_write_write                     : in  std_logic                     := 'X';             -- write
			sgdma_rx_m_write_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			sgdma_tx_m_read_address                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_tx_m_read_waitrequest                : out std_logic;                                        -- waitrequest
			sgdma_tx_m_read_read                       : in  std_logic                     := 'X';             -- read
			sgdma_tx_m_read_readdata                   : out std_logic_vector(31 downto 0);                    -- readdata
			sgdma_tx_m_read_readdatavalid              : out std_logic;                                        -- readdatavalid
			sgdma_bridge_s0_address                    : out std_logic_vector(30 downto 0);                    -- address
			sgdma_bridge_s0_write                      : out std_logic;                                        -- write
			sgdma_bridge_s0_read                       : out std_logic;                                        -- read
			sgdma_bridge_s0_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sgdma_bridge_s0_writedata                  : out std_logic_vector(31 downto 0);                    -- writedata
			sgdma_bridge_s0_burstcount                 : out std_logic_vector(0 downto 0);                     -- burstcount
			sgdma_bridge_s0_byteenable                 : out std_logic_vector(3 downto 0);                     -- byteenable
			sgdma_bridge_s0_readdatavalid              : in  std_logic                     := 'X';             -- readdatavalid
			sgdma_bridge_s0_waitrequest                : in  std_logic                     := 'X';             -- waitrequest
			sgdma_bridge_s0_debugaccess                : out std_logic                                         -- debugaccess
		);
	end component eth_std_main_system_ethernet_subsystem_mm_interconnect_2;

	component eth_std_main_system_ethernet_subsystem_avalon_st_adapter is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk        : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset      : in  std_logic                     := 'X';             -- reset
			in_0_data           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_0_valid          : in  std_logic                     := 'X';             -- valid
			in_0_ready          : out std_logic;                                        -- ready
			in_0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			in_0_empty          : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			in_0_error          : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- error
			out_0_data          : out std_logic_vector(31 downto 0);                    -- data
			out_0_valid         : out std_logic;                                        -- valid
			out_0_ready         : in  std_logic                     := 'X';             -- ready
			out_0_startofpacket : out std_logic;                                        -- startofpacket
			out_0_endofpacket   : out std_logic;                                        -- endofpacket
			out_0_empty         : out std_logic_vector(1 downto 0);                     -- empty
			out_0_error         : out std_logic_vector(5 downto 0)                      -- error
		);
	end component eth_std_main_system_ethernet_subsystem_avalon_st_adapter;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	component eth_std_main_system_ethernet_subsystem_ethernet_bridge is
		generic (
			DATA_WIDTH        : integer := 32;
			SYMBOL_WIDTH      : integer := 8;
			HDL_ADDR_WIDTH    : integer := 10;
			BURSTCOUNT_WIDTH  : integer := 1;
			PIPELINE_COMMAND  : integer := 1;
			PIPELINE_RESPONSE : integer := 1
		);
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset            : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(10 downto 0) := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(10 downto 0);                    -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic;                                        -- debugaccess
			s0_response      : out std_logic_vector(1 downto 0);                     -- response
			m0_response      : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- response
		);
	end component eth_std_main_system_ethernet_subsystem_ethernet_bridge;

	component eth_std_main_system_ethernet_subsystem_sgdma_bridge is
		generic (
			DATA_WIDTH        : integer := 32;
			SYMBOL_WIDTH      : integer := 8;
			HDL_ADDR_WIDTH    : integer := 10;
			BURSTCOUNT_WIDTH  : integer := 1;
			PIPELINE_COMMAND  : integer := 1;
			PIPELINE_RESPONSE : integer := 1
		);
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset            : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(30 downto 0) := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(30 downto 0);                    -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic;                                        -- debugaccess
			s0_response      : out std_logic_vector(1 downto 0);                     -- response
			m0_response      : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- response
		);
	end component eth_std_main_system_ethernet_subsystem_sgdma_bridge;

	signal sgdma_tx_out_valid                                 : std_logic;                     -- sgdma_tx:out_valid -> tse_mac:ff_tx_wren
	signal sgdma_tx_out_data                                  : std_logic_vector(31 downto 0); -- sgdma_tx:out_data -> tse_mac:ff_tx_data
	signal sgdma_tx_out_ready                                 : std_logic;                     -- tse_mac:ff_tx_rdy -> sgdma_tx:out_ready
	signal sgdma_tx_out_startofpacket                         : std_logic;                     -- sgdma_tx:out_startofpacket -> tse_mac:ff_tx_sop
	signal sgdma_tx_out_endofpacket                           : std_logic;                     -- sgdma_tx:out_endofpacket -> tse_mac:ff_tx_eop
	signal sgdma_tx_out_error                                 : std_logic;                     -- sgdma_tx:out_error -> tse_mac:ff_tx_err
	signal sgdma_tx_out_empty                                 : std_logic_vector(1 downto 0);  -- sgdma_tx:out_empty -> tse_mac:ff_tx_mod
	signal sgdma_tx_descriptor_read_readdata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:sgdma_tx_descriptor_read_readdata -> sgdma_tx:descriptor_read_readdata
	signal sgdma_tx_descriptor_read_waitrequest               : std_logic;                     -- mm_interconnect_0:sgdma_tx_descriptor_read_waitrequest -> sgdma_tx:descriptor_read_waitrequest
	signal sgdma_tx_descriptor_read_address                   : std_logic_vector(31 downto 0); -- sgdma_tx:descriptor_read_address -> mm_interconnect_0:sgdma_tx_descriptor_read_address
	signal sgdma_tx_descriptor_read_read                      : std_logic;                     -- sgdma_tx:descriptor_read_read -> mm_interconnect_0:sgdma_tx_descriptor_read_read
	signal sgdma_tx_descriptor_read_readdatavalid             : std_logic;                     -- mm_interconnect_0:sgdma_tx_descriptor_read_readdatavalid -> sgdma_tx:descriptor_read_readdatavalid
	signal sgdma_rx_descriptor_read_readdata                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:sgdma_rx_descriptor_read_readdata -> sgdma_rx:descriptor_read_readdata
	signal sgdma_rx_descriptor_read_waitrequest               : std_logic;                     -- mm_interconnect_0:sgdma_rx_descriptor_read_waitrequest -> sgdma_rx:descriptor_read_waitrequest
	signal sgdma_rx_descriptor_read_address                   : std_logic_vector(31 downto 0); -- sgdma_rx:descriptor_read_address -> mm_interconnect_0:sgdma_rx_descriptor_read_address
	signal sgdma_rx_descriptor_read_read                      : std_logic;                     -- sgdma_rx:descriptor_read_read -> mm_interconnect_0:sgdma_rx_descriptor_read_read
	signal sgdma_rx_descriptor_read_readdatavalid             : std_logic;                     -- mm_interconnect_0:sgdma_rx_descriptor_read_readdatavalid -> sgdma_rx:descriptor_read_readdatavalid
	signal sgdma_tx_descriptor_write_waitrequest              : std_logic;                     -- mm_interconnect_0:sgdma_tx_descriptor_write_waitrequest -> sgdma_tx:descriptor_write_waitrequest
	signal sgdma_tx_descriptor_write_address                  : std_logic_vector(31 downto 0); -- sgdma_tx:descriptor_write_address -> mm_interconnect_0:sgdma_tx_descriptor_write_address
	signal sgdma_tx_descriptor_write_write                    : std_logic;                     -- sgdma_tx:descriptor_write_write -> mm_interconnect_0:sgdma_tx_descriptor_write_write
	signal sgdma_tx_descriptor_write_writedata                : std_logic_vector(31 downto 0); -- sgdma_tx:descriptor_write_writedata -> mm_interconnect_0:sgdma_tx_descriptor_write_writedata
	signal sgdma_rx_descriptor_write_waitrequest              : std_logic;                     -- mm_interconnect_0:sgdma_rx_descriptor_write_waitrequest -> sgdma_rx:descriptor_write_waitrequest
	signal sgdma_rx_descriptor_write_address                  : std_logic_vector(31 downto 0); -- sgdma_rx:descriptor_write_address -> mm_interconnect_0:sgdma_rx_descriptor_write_address
	signal sgdma_rx_descriptor_write_write                    : std_logic;                     -- sgdma_rx:descriptor_write_write -> mm_interconnect_0:sgdma_rx_descriptor_write_write
	signal sgdma_rx_descriptor_write_writedata                : std_logic_vector(31 downto 0); -- sgdma_rx:descriptor_write_writedata -> mm_interconnect_0:sgdma_rx_descriptor_write_writedata
	signal mm_interconnect_0_descriptor_memory_s1_chipselect  : std_logic;                     -- mm_interconnect_0:descriptor_memory_s1_chipselect -> descriptor_memory:chipselect
	signal mm_interconnect_0_descriptor_memory_s1_readdata    : std_logic_vector(31 downto 0); -- descriptor_memory:readdata -> mm_interconnect_0:descriptor_memory_s1_readdata
	signal mm_interconnect_0_descriptor_memory_s1_address     : std_logic_vector(10 downto 0); -- mm_interconnect_0:descriptor_memory_s1_address -> descriptor_memory:address
	signal mm_interconnect_0_descriptor_memory_s1_byteenable  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:descriptor_memory_s1_byteenable -> descriptor_memory:byteenable
	signal mm_interconnect_0_descriptor_memory_s1_write       : std_logic;                     -- mm_interconnect_0:descriptor_memory_s1_write -> descriptor_memory:write
	signal mm_interconnect_0_descriptor_memory_s1_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_0:descriptor_memory_s1_writedata -> descriptor_memory:writedata
	signal mm_interconnect_0_descriptor_memory_s1_clken       : std_logic;                     -- mm_interconnect_0:descriptor_memory_s1_clken -> descriptor_memory:clken
	signal ethernet_bridge_m0_waitrequest                     : std_logic;                     -- mm_interconnect_1:ethernet_bridge_m0_waitrequest -> ethernet_bridge:m0_waitrequest
	signal ethernet_bridge_m0_readdata                        : std_logic_vector(31 downto 0); -- mm_interconnect_1:ethernet_bridge_m0_readdata -> ethernet_bridge:m0_readdata
	signal ethernet_bridge_m0_debugaccess                     : std_logic;                     -- ethernet_bridge:m0_debugaccess -> mm_interconnect_1:ethernet_bridge_m0_debugaccess
	signal ethernet_bridge_m0_address                         : std_logic_vector(10 downto 0); -- ethernet_bridge:m0_address -> mm_interconnect_1:ethernet_bridge_m0_address
	signal ethernet_bridge_m0_read                            : std_logic;                     -- ethernet_bridge:m0_read -> mm_interconnect_1:ethernet_bridge_m0_read
	signal ethernet_bridge_m0_byteenable                      : std_logic_vector(3 downto 0);  -- ethernet_bridge:m0_byteenable -> mm_interconnect_1:ethernet_bridge_m0_byteenable
	signal ethernet_bridge_m0_readdatavalid                   : std_logic;                     -- mm_interconnect_1:ethernet_bridge_m0_readdatavalid -> ethernet_bridge:m0_readdatavalid
	signal ethernet_bridge_m0_writedata                       : std_logic_vector(31 downto 0); -- ethernet_bridge:m0_writedata -> mm_interconnect_1:ethernet_bridge_m0_writedata
	signal ethernet_bridge_m0_write                           : std_logic;                     -- ethernet_bridge:m0_write -> mm_interconnect_1:ethernet_bridge_m0_write
	signal ethernet_bridge_m0_burstcount                      : std_logic_vector(0 downto 0);  -- ethernet_bridge:m0_burstcount -> mm_interconnect_1:ethernet_bridge_m0_burstcount
	signal mm_interconnect_1_tse_mac_control_port_readdata    : std_logic_vector(31 downto 0); -- tse_mac:reg_data_out -> mm_interconnect_1:tse_mac_control_port_readdata
	signal mm_interconnect_1_tse_mac_control_port_waitrequest : std_logic;                     -- tse_mac:reg_busy -> mm_interconnect_1:tse_mac_control_port_waitrequest
	signal mm_interconnect_1_tse_mac_control_port_address     : std_logic_vector(7 downto 0);  -- mm_interconnect_1:tse_mac_control_port_address -> tse_mac:reg_addr
	signal mm_interconnect_1_tse_mac_control_port_read        : std_logic;                     -- mm_interconnect_1:tse_mac_control_port_read -> tse_mac:reg_rd
	signal mm_interconnect_1_tse_mac_control_port_write       : std_logic;                     -- mm_interconnect_1:tse_mac_control_port_write -> tse_mac:reg_wr
	signal mm_interconnect_1_tse_mac_control_port_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_1:tse_mac_control_port_writedata -> tse_mac:reg_data_in
	signal mm_interconnect_1_sgdma_tx_csr_chipselect          : std_logic;                     -- mm_interconnect_1:sgdma_tx_csr_chipselect -> sgdma_tx:csr_chipselect
	signal mm_interconnect_1_sgdma_tx_csr_readdata            : std_logic_vector(31 downto 0); -- sgdma_tx:csr_readdata -> mm_interconnect_1:sgdma_tx_csr_readdata
	signal mm_interconnect_1_sgdma_tx_csr_address             : std_logic_vector(3 downto 0);  -- mm_interconnect_1:sgdma_tx_csr_address -> sgdma_tx:csr_address
	signal mm_interconnect_1_sgdma_tx_csr_read                : std_logic;                     -- mm_interconnect_1:sgdma_tx_csr_read -> sgdma_tx:csr_read
	signal mm_interconnect_1_sgdma_tx_csr_write               : std_logic;                     -- mm_interconnect_1:sgdma_tx_csr_write -> sgdma_tx:csr_write
	signal mm_interconnect_1_sgdma_tx_csr_writedata           : std_logic_vector(31 downto 0); -- mm_interconnect_1:sgdma_tx_csr_writedata -> sgdma_tx:csr_writedata
	signal mm_interconnect_1_sgdma_rx_csr_chipselect          : std_logic;                     -- mm_interconnect_1:sgdma_rx_csr_chipselect -> sgdma_rx:csr_chipselect
	signal mm_interconnect_1_sgdma_rx_csr_readdata            : std_logic_vector(31 downto 0); -- sgdma_rx:csr_readdata -> mm_interconnect_1:sgdma_rx_csr_readdata
	signal mm_interconnect_1_sgdma_rx_csr_address             : std_logic_vector(3 downto 0);  -- mm_interconnect_1:sgdma_rx_csr_address -> sgdma_rx:csr_address
	signal mm_interconnect_1_sgdma_rx_csr_read                : std_logic;                     -- mm_interconnect_1:sgdma_rx_csr_read -> sgdma_rx:csr_read
	signal mm_interconnect_1_sgdma_rx_csr_write               : std_logic;                     -- mm_interconnect_1:sgdma_rx_csr_write -> sgdma_rx:csr_write
	signal mm_interconnect_1_sgdma_rx_csr_writedata           : std_logic_vector(31 downto 0); -- mm_interconnect_1:sgdma_rx_csr_writedata -> sgdma_rx:csr_writedata
	signal sgdma_tx_m_read_readdata                           : std_logic_vector(31 downto 0); -- mm_interconnect_2:sgdma_tx_m_read_readdata -> sgdma_tx:m_read_readdata
	signal sgdma_tx_m_read_waitrequest                        : std_logic;                     -- mm_interconnect_2:sgdma_tx_m_read_waitrequest -> sgdma_tx:m_read_waitrequest
	signal sgdma_tx_m_read_address                            : std_logic_vector(31 downto 0); -- sgdma_tx:m_read_address -> mm_interconnect_2:sgdma_tx_m_read_address
	signal sgdma_tx_m_read_read                               : std_logic;                     -- sgdma_tx:m_read_read -> mm_interconnect_2:sgdma_tx_m_read_read
	signal sgdma_tx_m_read_readdatavalid                      : std_logic;                     -- mm_interconnect_2:sgdma_tx_m_read_readdatavalid -> sgdma_tx:m_read_readdatavalid
	signal sgdma_rx_m_write_waitrequest                       : std_logic;                     -- mm_interconnect_2:sgdma_rx_m_write_waitrequest -> sgdma_rx:m_write_waitrequest
	signal sgdma_rx_m_write_address                           : std_logic_vector(31 downto 0); -- sgdma_rx:m_write_address -> mm_interconnect_2:sgdma_rx_m_write_address
	signal sgdma_rx_m_write_byteenable                        : std_logic_vector(3 downto 0);  -- sgdma_rx:m_write_byteenable -> mm_interconnect_2:sgdma_rx_m_write_byteenable
	signal sgdma_rx_m_write_write                             : std_logic;                     -- sgdma_rx:m_write_write -> mm_interconnect_2:sgdma_rx_m_write_write
	signal sgdma_rx_m_write_writedata                         : std_logic_vector(31 downto 0); -- sgdma_rx:m_write_writedata -> mm_interconnect_2:sgdma_rx_m_write_writedata
	signal mm_interconnect_2_sgdma_bridge_s0_readdata         : std_logic_vector(31 downto 0); -- sgdma_bridge:s0_readdata -> mm_interconnect_2:sgdma_bridge_s0_readdata
	signal mm_interconnect_2_sgdma_bridge_s0_waitrequest      : std_logic;                     -- sgdma_bridge:s0_waitrequest -> mm_interconnect_2:sgdma_bridge_s0_waitrequest
	signal mm_interconnect_2_sgdma_bridge_s0_debugaccess      : std_logic;                     -- mm_interconnect_2:sgdma_bridge_s0_debugaccess -> sgdma_bridge:s0_debugaccess
	signal mm_interconnect_2_sgdma_bridge_s0_address          : std_logic_vector(30 downto 0); -- mm_interconnect_2:sgdma_bridge_s0_address -> sgdma_bridge:s0_address
	signal mm_interconnect_2_sgdma_bridge_s0_read             : std_logic;                     -- mm_interconnect_2:sgdma_bridge_s0_read -> sgdma_bridge:s0_read
	signal mm_interconnect_2_sgdma_bridge_s0_byteenable       : std_logic_vector(3 downto 0);  -- mm_interconnect_2:sgdma_bridge_s0_byteenable -> sgdma_bridge:s0_byteenable
	signal mm_interconnect_2_sgdma_bridge_s0_readdatavalid    : std_logic;                     -- sgdma_bridge:s0_readdatavalid -> mm_interconnect_2:sgdma_bridge_s0_readdatavalid
	signal mm_interconnect_2_sgdma_bridge_s0_write            : std_logic;                     -- mm_interconnect_2:sgdma_bridge_s0_write -> sgdma_bridge:s0_write
	signal mm_interconnect_2_sgdma_bridge_s0_writedata        : std_logic_vector(31 downto 0); -- mm_interconnect_2:sgdma_bridge_s0_writedata -> sgdma_bridge:s0_writedata
	signal mm_interconnect_2_sgdma_bridge_s0_burstcount       : std_logic_vector(0 downto 0);  -- mm_interconnect_2:sgdma_bridge_s0_burstcount -> sgdma_bridge:s0_burstcount
	signal tse_mac_receive_valid                              : std_logic;                     -- tse_mac:ff_rx_dval -> avalon_st_adapter:in_0_valid
	signal tse_mac_receive_data                               : std_logic_vector(31 downto 0); -- tse_mac:ff_rx_data -> avalon_st_adapter:in_0_data
	signal tse_mac_receive_ready                              : std_logic;                     -- avalon_st_adapter:in_0_ready -> tse_mac:ff_rx_rdy
	signal tse_mac_receive_startofpacket                      : std_logic;                     -- tse_mac:ff_rx_sop -> avalon_st_adapter:in_0_startofpacket
	signal tse_mac_receive_endofpacket                        : std_logic;                     -- tse_mac:ff_rx_eop -> avalon_st_adapter:in_0_endofpacket
	signal tse_mac_receive_error                              : std_logic_vector(5 downto 0);  -- tse_mac:rx_err -> avalon_st_adapter:in_0_error
	signal tse_mac_receive_empty                              : std_logic_vector(1 downto 0);  -- tse_mac:ff_rx_mod -> avalon_st_adapter:in_0_empty
	signal avalon_st_adapter_out_0_valid                      : std_logic;                     -- avalon_st_adapter:out_0_valid -> sgdma_rx:in_valid
	signal avalon_st_adapter_out_0_data                       : std_logic_vector(31 downto 0); -- avalon_st_adapter:out_0_data -> sgdma_rx:in_data
	signal avalon_st_adapter_out_0_ready                      : std_logic;                     -- sgdma_rx:in_ready -> avalon_st_adapter:out_0_ready
	signal avalon_st_adapter_out_0_startofpacket              : std_logic;                     -- avalon_st_adapter:out_0_startofpacket -> sgdma_rx:in_startofpacket
	signal avalon_st_adapter_out_0_endofpacket                : std_logic;                     -- avalon_st_adapter:out_0_endofpacket -> sgdma_rx:in_endofpacket
	signal avalon_st_adapter_out_0_error                      : std_logic_vector(5 downto 0);  -- avalon_st_adapter:out_0_error -> sgdma_rx:in_error
	signal avalon_st_adapter_out_0_empty                      : std_logic_vector(1 downto 0);  -- avalon_st_adapter:out_0_empty -> sgdma_rx:in_empty
	signal rst_controller_reset_out_reset                     : std_logic;                     -- rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, descriptor_memory:reset, descriptor_memory:reset2, ethernet_bridge:reset, mm_interconnect_0:sgdma_tx_reset_reset_bridge_in_reset_reset, mm_interconnect_1:ethernet_bridge_reset_reset_bridge_in_reset_reset, mm_interconnect_2:sgdma_tx_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset, sgdma_bridge:reset, tse_mac:reset]
	signal rst_controller_reset_out_reset_req                 : std_logic;                     -- rst_controller:reset_req -> [descriptor_memory:reset_req, descriptor_memory:reset_req2, rst_translator:reset_req_in]
	signal ethernet_subsys_reset_in_reset_n_ports_inv         : std_logic;                     -- ethernet_subsys_reset_in_reset_n:inv -> rst_controller:reset_in0
	signal rst_controller_reset_out_reset_ports_inv           : std_logic;                     -- rst_controller_reset_out_reset:inv -> [sgdma_rx:system_reset_n, sgdma_tx:system_reset_n]

begin

	descriptor_memory : component eth_std_main_system_ethernet_subsystem_descriptor_memory
		port map (
			clk         => ethernet_subsys_clk_in_clk,                        --   clk1.clk
			address     => mm_interconnect_0_descriptor_memory_s1_address,    --     s1.address
			clken       => mm_interconnect_0_descriptor_memory_s1_clken,      --       .clken
			chipselect  => mm_interconnect_0_descriptor_memory_s1_chipselect, --       .chipselect
			write       => mm_interconnect_0_descriptor_memory_s1_write,      --       .write
			readdata    => mm_interconnect_0_descriptor_memory_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_0_descriptor_memory_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_0_descriptor_memory_s1_byteenable, --       .byteenable
			reset       => rst_controller_reset_out_reset,                    -- reset1.reset
			reset_req   => rst_controller_reset_out_reset_req,                --       .reset_req
			address2    => descriptor_memory_s2_address,                      --     s2.address
			chipselect2 => descriptor_memory_s2_chipselect,                   --       .chipselect
			clken2      => descriptor_memory_s2_clken,                        --       .clken
			write2      => descriptor_memory_s2_write,                        --       .write
			readdata2   => descriptor_memory_s2_readdata,                     --       .readdata
			writedata2  => descriptor_memory_s2_writedata,                    --       .writedata
			byteenable2 => descriptor_memory_s2_byteenable,                   --       .byteenable
			clk2        => ethernet_subsys_clk_in_clk,                        --   clk2.clk
			reset2      => rst_controller_reset_out_reset,                    -- reset2.reset
			reset_req2  => rst_controller_reset_out_reset_req,                --       .reset_req
			freeze      => '0'                                                -- (terminated)
		);

	ethernet_bridge : component eth_std_main_system_ethernet_subsystem_ethernet_bridge
		generic map (
			DATA_WIDTH        => 32,
			SYMBOL_WIDTH      => 8,
			HDL_ADDR_WIDTH    => 11,
			BURSTCOUNT_WIDTH  => 1,
			PIPELINE_COMMAND  => 1,
			PIPELINE_RESPONSE => 1
		)
		port map (
			clk              => ethernet_subsys_clk_in_clk,       --   clk.clk
			reset            => rst_controller_reset_out_reset,   -- reset.reset
			s0_waitrequest   => ethernet_bridge_s0_waitrequest,   --    s0.waitrequest
			s0_readdata      => ethernet_bridge_s0_readdata,      --      .readdata
			s0_readdatavalid => ethernet_bridge_s0_readdatavalid, --      .readdatavalid
			s0_burstcount    => ethernet_bridge_s0_burstcount,    --      .burstcount
			s0_writedata     => ethernet_bridge_s0_writedata,     --      .writedata
			s0_address       => ethernet_bridge_s0_address,       --      .address
			s0_write         => ethernet_bridge_s0_write,         --      .write
			s0_read          => ethernet_bridge_s0_read,          --      .read
			s0_byteenable    => ethernet_bridge_s0_byteenable,    --      .byteenable
			s0_debugaccess   => ethernet_bridge_s0_debugaccess,   --      .debugaccess
			m0_waitrequest   => ethernet_bridge_m0_waitrequest,   --    m0.waitrequest
			m0_readdata      => ethernet_bridge_m0_readdata,      --      .readdata
			m0_readdatavalid => ethernet_bridge_m0_readdatavalid, --      .readdatavalid
			m0_burstcount    => ethernet_bridge_m0_burstcount,    --      .burstcount
			m0_writedata     => ethernet_bridge_m0_writedata,     --      .writedata
			m0_address       => ethernet_bridge_m0_address,       --      .address
			m0_write         => ethernet_bridge_m0_write,         --      .write
			m0_read          => ethernet_bridge_m0_read,          --      .read
			m0_byteenable    => ethernet_bridge_m0_byteenable,    --      .byteenable
			m0_debugaccess   => ethernet_bridge_m0_debugaccess,   --      .debugaccess
			s0_response      => open,                             -- (terminated)
			m0_response      => "00"                              -- (terminated)
		);

	sgdma_bridge : component eth_std_main_system_ethernet_subsystem_sgdma_bridge
		generic map (
			DATA_WIDTH        => 32,
			SYMBOL_WIDTH      => 8,
			HDL_ADDR_WIDTH    => 31,
			BURSTCOUNT_WIDTH  => 1,
			PIPELINE_COMMAND  => 1,
			PIPELINE_RESPONSE => 1
		)
		port map (
			clk              => ethernet_subsys_clk_in_clk,                      --   clk.clk
			reset            => rst_controller_reset_out_reset,                  -- reset.reset
			s0_waitrequest   => mm_interconnect_2_sgdma_bridge_s0_waitrequest,   --    s0.waitrequest
			s0_readdata      => mm_interconnect_2_sgdma_bridge_s0_readdata,      --      .readdata
			s0_readdatavalid => mm_interconnect_2_sgdma_bridge_s0_readdatavalid, --      .readdatavalid
			s0_burstcount    => mm_interconnect_2_sgdma_bridge_s0_burstcount,    --      .burstcount
			s0_writedata     => mm_interconnect_2_sgdma_bridge_s0_writedata,     --      .writedata
			s0_address       => mm_interconnect_2_sgdma_bridge_s0_address,       --      .address
			s0_write         => mm_interconnect_2_sgdma_bridge_s0_write,         --      .write
			s0_read          => mm_interconnect_2_sgdma_bridge_s0_read,          --      .read
			s0_byteenable    => mm_interconnect_2_sgdma_bridge_s0_byteenable,    --      .byteenable
			s0_debugaccess   => mm_interconnect_2_sgdma_bridge_s0_debugaccess,   --      .debugaccess
			m0_waitrequest   => sgdma_bridge_m0_waitrequest,                     --    m0.waitrequest
			m0_readdata      => sgdma_bridge_m0_readdata,                        --      .readdata
			m0_readdatavalid => sgdma_bridge_m0_readdatavalid,                   --      .readdatavalid
			m0_burstcount    => sgdma_bridge_m0_burstcount,                      --      .burstcount
			m0_writedata     => sgdma_bridge_m0_writedata,                       --      .writedata
			m0_address       => sgdma_bridge_m0_address,                         --      .address
			m0_write         => sgdma_bridge_m0_write,                           --      .write
			m0_read          => sgdma_bridge_m0_read,                            --      .read
			m0_byteenable    => sgdma_bridge_m0_byteenable,                      --      .byteenable
			m0_debugaccess   => sgdma_bridge_m0_debugaccess,                     --      .debugaccess
			s0_response      => open,                                            -- (terminated)
			m0_response      => "00"                                             -- (terminated)
		);

	sgdma_rx : component eth_std_main_system_ethernet_subsystem_sgdma_rx
		port map (
			clk                           => ethernet_subsys_clk_in_clk,                --              clk.clk
			system_reset_n                => rst_controller_reset_out_reset_ports_inv,  --            reset.reset_n
			csr_chipselect                => mm_interconnect_1_sgdma_rx_csr_chipselect, --              csr.chipselect
			csr_address                   => mm_interconnect_1_sgdma_rx_csr_address,    --                 .address
			csr_read                      => mm_interconnect_1_sgdma_rx_csr_read,       --                 .read
			csr_write                     => mm_interconnect_1_sgdma_rx_csr_write,      --                 .write
			csr_writedata                 => mm_interconnect_1_sgdma_rx_csr_writedata,  --                 .writedata
			csr_readdata                  => mm_interconnect_1_sgdma_rx_csr_readdata,   --                 .readdata
			descriptor_read_readdata      => sgdma_rx_descriptor_read_readdata,         --  descriptor_read.readdata
			descriptor_read_readdatavalid => sgdma_rx_descriptor_read_readdatavalid,    --                 .readdatavalid
			descriptor_read_waitrequest   => sgdma_rx_descriptor_read_waitrequest,      --                 .waitrequest
			descriptor_read_address       => sgdma_rx_descriptor_read_address,          --                 .address
			descriptor_read_read          => sgdma_rx_descriptor_read_read,             --                 .read
			descriptor_write_waitrequest  => sgdma_rx_descriptor_write_waitrequest,     -- descriptor_write.waitrequest
			descriptor_write_address      => sgdma_rx_descriptor_write_address,         --                 .address
			descriptor_write_write        => sgdma_rx_descriptor_write_write,           --                 .write
			descriptor_write_writedata    => sgdma_rx_descriptor_write_writedata,       --                 .writedata
			csr_irq                       => sgdma_rx_csr_irq_irq,                      --          csr_irq.irq
			in_startofpacket              => avalon_st_adapter_out_0_startofpacket,     --               in.startofpacket
			in_endofpacket                => avalon_st_adapter_out_0_endofpacket,       --                 .endofpacket
			in_data                       => avalon_st_adapter_out_0_data,              --                 .data
			in_valid                      => avalon_st_adapter_out_0_valid,             --                 .valid
			in_ready                      => avalon_st_adapter_out_0_ready,             --                 .ready
			in_empty                      => avalon_st_adapter_out_0_empty,             --                 .empty
			in_error                      => avalon_st_adapter_out_0_error,             --                 .error
			m_write_waitrequest           => sgdma_rx_m_write_waitrequest,              --          m_write.waitrequest
			m_write_address               => sgdma_rx_m_write_address,                  --                 .address
			m_write_write                 => sgdma_rx_m_write_write,                    --                 .write
			m_write_writedata             => sgdma_rx_m_write_writedata,                --                 .writedata
			m_write_byteenable            => sgdma_rx_m_write_byteenable                --                 .byteenable
		);

	sgdma_tx : component eth_std_main_system_ethernet_subsystem_sgdma_tx
		port map (
			clk                           => ethernet_subsys_clk_in_clk,                --              clk.clk
			system_reset_n                => rst_controller_reset_out_reset_ports_inv,  --            reset.reset_n
			csr_chipselect                => mm_interconnect_1_sgdma_tx_csr_chipselect, --              csr.chipselect
			csr_address                   => mm_interconnect_1_sgdma_tx_csr_address,    --                 .address
			csr_read                      => mm_interconnect_1_sgdma_tx_csr_read,       --                 .read
			csr_write                     => mm_interconnect_1_sgdma_tx_csr_write,      --                 .write
			csr_writedata                 => mm_interconnect_1_sgdma_tx_csr_writedata,  --                 .writedata
			csr_readdata                  => mm_interconnect_1_sgdma_tx_csr_readdata,   --                 .readdata
			descriptor_read_readdata      => sgdma_tx_descriptor_read_readdata,         --  descriptor_read.readdata
			descriptor_read_readdatavalid => sgdma_tx_descriptor_read_readdatavalid,    --                 .readdatavalid
			descriptor_read_waitrequest   => sgdma_tx_descriptor_read_waitrequest,      --                 .waitrequest
			descriptor_read_address       => sgdma_tx_descriptor_read_address,          --                 .address
			descriptor_read_read          => sgdma_tx_descriptor_read_read,             --                 .read
			descriptor_write_waitrequest  => sgdma_tx_descriptor_write_waitrequest,     -- descriptor_write.waitrequest
			descriptor_write_address      => sgdma_tx_descriptor_write_address,         --                 .address
			descriptor_write_write        => sgdma_tx_descriptor_write_write,           --                 .write
			descriptor_write_writedata    => sgdma_tx_descriptor_write_writedata,       --                 .writedata
			csr_irq                       => sgdma_tx_csr_irq_irq,                      --          csr_irq.irq
			m_read_readdata               => sgdma_tx_m_read_readdata,                  --           m_read.readdata
			m_read_readdatavalid          => sgdma_tx_m_read_readdatavalid,             --                 .readdatavalid
			m_read_waitrequest            => sgdma_tx_m_read_waitrequest,               --                 .waitrequest
			m_read_address                => sgdma_tx_m_read_address,                   --                 .address
			m_read_read                   => sgdma_tx_m_read_read,                      --                 .read
			out_data                      => sgdma_tx_out_data,                         --              out.data
			out_valid                     => sgdma_tx_out_valid,                        --                 .valid
			out_ready                     => sgdma_tx_out_ready,                        --                 .ready
			out_endofpacket               => sgdma_tx_out_endofpacket,                  --                 .endofpacket
			out_startofpacket             => sgdma_tx_out_startofpacket,                --                 .startofpacket
			out_empty                     => sgdma_tx_out_empty,                        --                 .empty
			out_error                     => sgdma_tx_out_error                         --                 .error
		);

	tse_mac : component eth_std_main_system_ethernet_subsystem_tse_mac
		port map (
			clk           => ethernet_subsys_clk_in_clk,                         -- control_port_clock_connection.clk
			reset         => rst_controller_reset_out_reset,                     --              reset_connection.reset
			reg_addr      => mm_interconnect_1_tse_mac_control_port_address,     --                  control_port.address
			reg_data_out  => mm_interconnect_1_tse_mac_control_port_readdata,    --                              .readdata
			reg_rd        => mm_interconnect_1_tse_mac_control_port_read,        --                              .read
			reg_data_in   => mm_interconnect_1_tse_mac_control_port_writedata,   --                              .writedata
			reg_wr        => mm_interconnect_1_tse_mac_control_port_write,       --                              .write
			reg_busy      => mm_interconnect_1_tse_mac_control_port_waitrequest, --                              .waitrequest
			tx_clk        => tx_clock_clk,                                       --   pcs_mac_tx_clock_connection.clk
			rx_clk        => rx_clock_clk,                                       --   pcs_mac_rx_clock_connection.clk
			set_10        => mac_status_connection_set_10,                       --         mac_status_connection.set_10
			set_1000      => mac_status_connection_set_1000,                     --                              .set_1000
			eth_mode      => mac_status_connection_eth_mode,                     --                              .eth_mode
			ena_10        => mac_status_connection_ena_10,                       --                              .ena_10
			gm_rx_d       => mac_gmii_connection_gmii_rx_d,                      --           mac_gmii_connection.gmii_rx_d
			gm_rx_dv      => mac_gmii_connection_gmii_rx_dv,                     --                              .gmii_rx_dv
			gm_rx_err     => mac_gmii_connection_gmii_rx_err,                    --                              .gmii_rx_err
			gm_tx_d       => mac_gmii_connection_gmii_tx_d,                      --                              .gmii_tx_d
			gm_tx_en      => mac_gmii_connection_gmii_tx_en,                     --                              .gmii_tx_en
			gm_tx_err     => mac_gmii_connection_gmii_tx_err,                    --                              .gmii_tx_err
			m_rx_d        => mac_mii_connection_mii_rx_d,                        --            mac_mii_connection.mii_rx_d
			m_rx_en       => mac_mii_connection_mii_rx_dv,                       --                              .mii_rx_dv
			m_rx_err      => mac_mii_connection_mii_rx_err,                      --                              .mii_rx_err
			m_tx_d        => mac_mii_connection_mii_tx_d,                        --                              .mii_tx_d
			m_tx_en       => mac_mii_connection_mii_tx_en,                       --                              .mii_tx_en
			m_tx_err      => mac_mii_connection_mii_tx_err,                      --                              .mii_tx_err
			m_rx_crs      => mac_mii_connection_mii_crs,                         --                              .mii_crs
			m_rx_col      => mac_mii_connection_mii_col,                         --                              .mii_col
			ff_rx_clk     => ethernet_subsys_clk_in_clk,                         --      receive_clock_connection.clk
			ff_tx_clk     => ethernet_subsys_clk_in_clk,                         --     transmit_clock_connection.clk
			ff_rx_data    => tse_mac_receive_data,                               --                       receive.data
			ff_rx_eop     => tse_mac_receive_endofpacket,                        --                              .endofpacket
			rx_err        => tse_mac_receive_error,                              --                              .error
			ff_rx_mod     => tse_mac_receive_empty,                              --                              .empty
			ff_rx_rdy     => tse_mac_receive_ready,                              --                              .ready
			ff_rx_sop     => tse_mac_receive_startofpacket,                      --                              .startofpacket
			ff_rx_dval    => tse_mac_receive_valid,                              --                              .valid
			ff_tx_data    => sgdma_tx_out_data,                                  --                      transmit.data
			ff_tx_eop     => sgdma_tx_out_endofpacket,                           --                              .endofpacket
			ff_tx_err     => sgdma_tx_out_error,                                 --                              .error
			ff_tx_mod     => sgdma_tx_out_empty,                                 --                              .empty
			ff_tx_rdy     => sgdma_tx_out_ready,                                 --                              .ready
			ff_tx_sop     => sgdma_tx_out_startofpacket,                         --                              .startofpacket
			ff_tx_wren    => sgdma_tx_out_valid,                                 --                              .valid
			mdc           => mac_mdio_connection_mdc,                            --           mac_mdio_connection.mdc
			mdio_in       => mac_mdio_connection_mdio_in,                        --                              .mdio_in
			mdio_out      => mac_mdio_connection_mdio_out,                       --                              .mdio_out
			mdio_oen      => mac_mdio_connection_mdio_oen,                       --                              .mdio_oen
			xon_gen       => misc_connection_xon_gen,                            --           mac_misc_connection.xon_gen
			xoff_gen      => misc_connection_xoff_gen,                           --                              .xoff_gen
			ff_tx_crc_fwd => misc_connection_ff_tx_crc_fwd,                      --                              .ff_tx_crc_fwd
			ff_tx_septy   => misc_connection_ff_tx_septy,                        --                              .ff_tx_septy
			tx_ff_uflow   => misc_connection_tx_ff_uflow,                        --                              .tx_ff_uflow
			ff_tx_a_full  => misc_connection_ff_tx_a_full,                       --                              .ff_tx_a_full
			ff_tx_a_empty => misc_connection_ff_tx_a_empty,                      --                              .ff_tx_a_empty
			rx_err_stat   => misc_connection_rx_err_stat,                        --                              .rx_err_stat
			rx_frm_type   => misc_connection_rx_frm_type,                        --                              .rx_frm_type
			ff_rx_dsav    => misc_connection_ff_rx_dsav,                         --                              .ff_rx_dsav
			ff_rx_a_full  => misc_connection_ff_rx_a_full,                       --                              .ff_rx_a_full
			ff_rx_a_empty => misc_connection_ff_rx_a_empty                       --                              .ff_rx_a_empty
		);

	mm_interconnect_0 : component eth_std_main_system_ethernet_subsystem_mm_interconnect_0
		port map (
			clk_clk_clk                                => ethernet_subsys_clk_in_clk,                        --                              clk_clk.clk
			sgdma_tx_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                    -- sgdma_tx_reset_reset_bridge_in_reset.reset
			sgdma_rx_descriptor_read_address           => sgdma_rx_descriptor_read_address,                  --             sgdma_rx_descriptor_read.address
			sgdma_rx_descriptor_read_waitrequest       => sgdma_rx_descriptor_read_waitrequest,              --                                     .waitrequest
			sgdma_rx_descriptor_read_read              => sgdma_rx_descriptor_read_read,                     --                                     .read
			sgdma_rx_descriptor_read_readdata          => sgdma_rx_descriptor_read_readdata,                 --                                     .readdata
			sgdma_rx_descriptor_read_readdatavalid     => sgdma_rx_descriptor_read_readdatavalid,            --                                     .readdatavalid
			sgdma_rx_descriptor_write_address          => sgdma_rx_descriptor_write_address,                 --            sgdma_rx_descriptor_write.address
			sgdma_rx_descriptor_write_waitrequest      => sgdma_rx_descriptor_write_waitrequest,             --                                     .waitrequest
			sgdma_rx_descriptor_write_write            => sgdma_rx_descriptor_write_write,                   --                                     .write
			sgdma_rx_descriptor_write_writedata        => sgdma_rx_descriptor_write_writedata,               --                                     .writedata
			sgdma_tx_descriptor_read_address           => sgdma_tx_descriptor_read_address,                  --             sgdma_tx_descriptor_read.address
			sgdma_tx_descriptor_read_waitrequest       => sgdma_tx_descriptor_read_waitrequest,              --                                     .waitrequest
			sgdma_tx_descriptor_read_read              => sgdma_tx_descriptor_read_read,                     --                                     .read
			sgdma_tx_descriptor_read_readdata          => sgdma_tx_descriptor_read_readdata,                 --                                     .readdata
			sgdma_tx_descriptor_read_readdatavalid     => sgdma_tx_descriptor_read_readdatavalid,            --                                     .readdatavalid
			sgdma_tx_descriptor_write_address          => sgdma_tx_descriptor_write_address,                 --            sgdma_tx_descriptor_write.address
			sgdma_tx_descriptor_write_waitrequest      => sgdma_tx_descriptor_write_waitrequest,             --                                     .waitrequest
			sgdma_tx_descriptor_write_write            => sgdma_tx_descriptor_write_write,                   --                                     .write
			sgdma_tx_descriptor_write_writedata        => sgdma_tx_descriptor_write_writedata,               --                                     .writedata
			descriptor_memory_s1_address               => mm_interconnect_0_descriptor_memory_s1_address,    --                 descriptor_memory_s1.address
			descriptor_memory_s1_write                 => mm_interconnect_0_descriptor_memory_s1_write,      --                                     .write
			descriptor_memory_s1_readdata              => mm_interconnect_0_descriptor_memory_s1_readdata,   --                                     .readdata
			descriptor_memory_s1_writedata             => mm_interconnect_0_descriptor_memory_s1_writedata,  --                                     .writedata
			descriptor_memory_s1_byteenable            => mm_interconnect_0_descriptor_memory_s1_byteenable, --                                     .byteenable
			descriptor_memory_s1_chipselect            => mm_interconnect_0_descriptor_memory_s1_chipselect, --                                     .chipselect
			descriptor_memory_s1_clken                 => mm_interconnect_0_descriptor_memory_s1_clken       --                                     .clken
		);

	mm_interconnect_1 : component eth_std_main_system_ethernet_subsystem_mm_interconnect_1
		port map (
			clk_clk_clk                                       => ethernet_subsys_clk_in_clk,                         --                                     clk_clk.clk
			ethernet_bridge_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                     -- ethernet_bridge_reset_reset_bridge_in_reset.reset
			ethernet_bridge_m0_address                        => ethernet_bridge_m0_address,                         --                          ethernet_bridge_m0.address
			ethernet_bridge_m0_waitrequest                    => ethernet_bridge_m0_waitrequest,                     --                                            .waitrequest
			ethernet_bridge_m0_burstcount                     => ethernet_bridge_m0_burstcount,                      --                                            .burstcount
			ethernet_bridge_m0_byteenable                     => ethernet_bridge_m0_byteenable,                      --                                            .byteenable
			ethernet_bridge_m0_read                           => ethernet_bridge_m0_read,                            --                                            .read
			ethernet_bridge_m0_readdata                       => ethernet_bridge_m0_readdata,                        --                                            .readdata
			ethernet_bridge_m0_readdatavalid                  => ethernet_bridge_m0_readdatavalid,                   --                                            .readdatavalid
			ethernet_bridge_m0_write                          => ethernet_bridge_m0_write,                           --                                            .write
			ethernet_bridge_m0_writedata                      => ethernet_bridge_m0_writedata,                       --                                            .writedata
			ethernet_bridge_m0_debugaccess                    => ethernet_bridge_m0_debugaccess,                     --                                            .debugaccess
			sgdma_rx_csr_address                              => mm_interconnect_1_sgdma_rx_csr_address,             --                                sgdma_rx_csr.address
			sgdma_rx_csr_write                                => mm_interconnect_1_sgdma_rx_csr_write,               --                                            .write
			sgdma_rx_csr_read                                 => mm_interconnect_1_sgdma_rx_csr_read,                --                                            .read
			sgdma_rx_csr_readdata                             => mm_interconnect_1_sgdma_rx_csr_readdata,            --                                            .readdata
			sgdma_rx_csr_writedata                            => mm_interconnect_1_sgdma_rx_csr_writedata,           --                                            .writedata
			sgdma_rx_csr_chipselect                           => mm_interconnect_1_sgdma_rx_csr_chipselect,          --                                            .chipselect
			sgdma_tx_csr_address                              => mm_interconnect_1_sgdma_tx_csr_address,             --                                sgdma_tx_csr.address
			sgdma_tx_csr_write                                => mm_interconnect_1_sgdma_tx_csr_write,               --                                            .write
			sgdma_tx_csr_read                                 => mm_interconnect_1_sgdma_tx_csr_read,                --                                            .read
			sgdma_tx_csr_readdata                             => mm_interconnect_1_sgdma_tx_csr_readdata,            --                                            .readdata
			sgdma_tx_csr_writedata                            => mm_interconnect_1_sgdma_tx_csr_writedata,           --                                            .writedata
			sgdma_tx_csr_chipselect                           => mm_interconnect_1_sgdma_tx_csr_chipselect,          --                                            .chipselect
			tse_mac_control_port_address                      => mm_interconnect_1_tse_mac_control_port_address,     --                        tse_mac_control_port.address
			tse_mac_control_port_write                        => mm_interconnect_1_tse_mac_control_port_write,       --                                            .write
			tse_mac_control_port_read                         => mm_interconnect_1_tse_mac_control_port_read,        --                                            .read
			tse_mac_control_port_readdata                     => mm_interconnect_1_tse_mac_control_port_readdata,    --                                            .readdata
			tse_mac_control_port_writedata                    => mm_interconnect_1_tse_mac_control_port_writedata,   --                                            .writedata
			tse_mac_control_port_waitrequest                  => mm_interconnect_1_tse_mac_control_port_waitrequest  --                                            .waitrequest
		);

	mm_interconnect_2 : component eth_std_main_system_ethernet_subsystem_mm_interconnect_2
		port map (
			clk_clk_clk                                => ethernet_subsys_clk_in_clk,                      --                              clk_clk.clk
			sgdma_tx_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                  -- sgdma_tx_reset_reset_bridge_in_reset.reset
			sgdma_rx_m_write_address                   => sgdma_rx_m_write_address,                        --                     sgdma_rx_m_write.address
			sgdma_rx_m_write_waitrequest               => sgdma_rx_m_write_waitrequest,                    --                                     .waitrequest
			sgdma_rx_m_write_byteenable                => sgdma_rx_m_write_byteenable,                     --                                     .byteenable
			sgdma_rx_m_write_write                     => sgdma_rx_m_write_write,                          --                                     .write
			sgdma_rx_m_write_writedata                 => sgdma_rx_m_write_writedata,                      --                                     .writedata
			sgdma_tx_m_read_address                    => sgdma_tx_m_read_address,                         --                      sgdma_tx_m_read.address
			sgdma_tx_m_read_waitrequest                => sgdma_tx_m_read_waitrequest,                     --                                     .waitrequest
			sgdma_tx_m_read_read                       => sgdma_tx_m_read_read,                            --                                     .read
			sgdma_tx_m_read_readdata                   => sgdma_tx_m_read_readdata,                        --                                     .readdata
			sgdma_tx_m_read_readdatavalid              => sgdma_tx_m_read_readdatavalid,                   --                                     .readdatavalid
			sgdma_bridge_s0_address                    => mm_interconnect_2_sgdma_bridge_s0_address,       --                      sgdma_bridge_s0.address
			sgdma_bridge_s0_write                      => mm_interconnect_2_sgdma_bridge_s0_write,         --                                     .write
			sgdma_bridge_s0_read                       => mm_interconnect_2_sgdma_bridge_s0_read,          --                                     .read
			sgdma_bridge_s0_readdata                   => mm_interconnect_2_sgdma_bridge_s0_readdata,      --                                     .readdata
			sgdma_bridge_s0_writedata                  => mm_interconnect_2_sgdma_bridge_s0_writedata,     --                                     .writedata
			sgdma_bridge_s0_burstcount                 => mm_interconnect_2_sgdma_bridge_s0_burstcount,    --                                     .burstcount
			sgdma_bridge_s0_byteenable                 => mm_interconnect_2_sgdma_bridge_s0_byteenable,    --                                     .byteenable
			sgdma_bridge_s0_readdatavalid              => mm_interconnect_2_sgdma_bridge_s0_readdatavalid, --                                     .readdatavalid
			sgdma_bridge_s0_waitrequest                => mm_interconnect_2_sgdma_bridge_s0_waitrequest,   --                                     .waitrequest
			sgdma_bridge_s0_debugaccess                => mm_interconnect_2_sgdma_bridge_s0_debugaccess    --                                     .debugaccess
		);

	avalon_st_adapter : component eth_std_main_system_ethernet_subsystem_avalon_st_adapter
		generic map (
			inBitsPerSymbol => 8,
			inUsePackets    => 1,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 6,
			inUseEmptyPort  => 1,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 2,
			outDataWidth    => 32,
			outChannelWidth => 0,
			outErrorWidth   => 6,
			outUseEmptyPort => 1,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk        => ethernet_subsys_clk_in_clk,            -- in_clk_0.clk
			in_rst_0_reset      => rst_controller_reset_out_reset,        -- in_rst_0.reset
			in_0_data           => tse_mac_receive_data,                  --     in_0.data
			in_0_valid          => tse_mac_receive_valid,                 --         .valid
			in_0_ready          => tse_mac_receive_ready,                 --         .ready
			in_0_startofpacket  => tse_mac_receive_startofpacket,         --         .startofpacket
			in_0_endofpacket    => tse_mac_receive_endofpacket,           --         .endofpacket
			in_0_empty          => tse_mac_receive_empty,                 --         .empty
			in_0_error          => tse_mac_receive_error,                 --         .error
			out_0_data          => avalon_st_adapter_out_0_data,          --    out_0.data
			out_0_valid         => avalon_st_adapter_out_0_valid,         --         .valid
			out_0_ready         => avalon_st_adapter_out_0_ready,         --         .ready
			out_0_startofpacket => avalon_st_adapter_out_0_startofpacket, --         .startofpacket
			out_0_endofpacket   => avalon_st_adapter_out_0_endofpacket,   --         .endofpacket
			out_0_empty         => avalon_st_adapter_out_0_empty,         --         .empty
			out_0_error         => avalon_st_adapter_out_0_error          --         .error
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => ethernet_subsys_reset_in_reset_n_ports_inv, -- reset_in0.reset
			clk            => ethernet_subsys_clk_in_clk,                 --       clk.clk
			reset_out      => rst_controller_reset_out_reset,             -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,         --          .reset_req
			reset_req_in0  => '0',                                        -- (terminated)
			reset_in1      => '0',                                        -- (terminated)
			reset_req_in1  => '0',                                        -- (terminated)
			reset_in2      => '0',                                        -- (terminated)
			reset_req_in2  => '0',                                        -- (terminated)
			reset_in3      => '0',                                        -- (terminated)
			reset_req_in3  => '0',                                        -- (terminated)
			reset_in4      => '0',                                        -- (terminated)
			reset_req_in4  => '0',                                        -- (terminated)
			reset_in5      => '0',                                        -- (terminated)
			reset_req_in5  => '0',                                        -- (terminated)
			reset_in6      => '0',                                        -- (terminated)
			reset_req_in6  => '0',                                        -- (terminated)
			reset_in7      => '0',                                        -- (terminated)
			reset_req_in7  => '0',                                        -- (terminated)
			reset_in8      => '0',                                        -- (terminated)
			reset_req_in8  => '0',                                        -- (terminated)
			reset_in9      => '0',                                        -- (terminated)
			reset_req_in9  => '0',                                        -- (terminated)
			reset_in10     => '0',                                        -- (terminated)
			reset_req_in10 => '0',                                        -- (terminated)
			reset_in11     => '0',                                        -- (terminated)
			reset_req_in11 => '0',                                        -- (terminated)
			reset_in12     => '0',                                        -- (terminated)
			reset_req_in12 => '0',                                        -- (terminated)
			reset_in13     => '0',                                        -- (terminated)
			reset_req_in13 => '0',                                        -- (terminated)
			reset_in14     => '0',                                        -- (terminated)
			reset_req_in14 => '0',                                        -- (terminated)
			reset_in15     => '0',                                        -- (terminated)
			reset_req_in15 => '0'                                         -- (terminated)
		);

	ethernet_subsys_reset_in_reset_n_ports_inv <= not ethernet_subsys_reset_in_reset_n;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of eth_std_main_system_ethernet_subsystem
