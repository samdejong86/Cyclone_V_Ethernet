-- peripheral_system.vhd

-- Generated using ACDS version 16.1 196

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity peripheral_system is
	port (
		button_pio_external_connection_export : in  std_logic_vector(2 downto 0)  := (others => '0'); -- button_pio_external_connection.export
		button_pio_irq_irq                    : out std_logic;                                        --                 button_pio_irq.irq
		high_res_timer_irq_irq                : out std_logic;                                        --             high_res_timer_irq.irq
		jtag_uart_irq_irq                     : out std_logic;                                        --                  jtag_uart_irq.irq
		led_pio_external_connection_export    : out std_logic_vector(7 downto 0);                     --    led_pio_external_connection.export
		peripheral_bridge_s0_waitrequest      : out std_logic;                                        --           peripheral_bridge_s0.waitrequest
		peripheral_bridge_s0_readdata         : out std_logic_vector(31 downto 0);                    --                               .readdata
		peripheral_bridge_s0_readdatavalid    : out std_logic;                                        --                               .readdatavalid
		peripheral_bridge_s0_burstcount       : in  std_logic_vector(0 downto 0)  := (others => '0'); --                               .burstcount
		peripheral_bridge_s0_writedata        : in  std_logic_vector(31 downto 0) := (others => '0'); --                               .writedata
		peripheral_bridge_s0_address          : in  std_logic_vector(7 downto 0)  := (others => '0'); --                               .address
		peripheral_bridge_s0_write            : in  std_logic                     := '0';             --                               .write
		peripheral_bridge_s0_read             : in  std_logic                     := '0';             --                               .read
		peripheral_bridge_s0_byteenable       : in  std_logic_vector(3 downto 0)  := (others => '0'); --                               .byteenable
		peripheral_bridge_s0_debugaccess      : in  std_logic                     := '0';             --                               .debugaccess
		peripheral_subsys_clk_in_clk          : in  std_logic                     := '0';             --       peripheral_subsys_clk_in.clk
		peripheral_subsys_reset_in_reset_n    : in  std_logic                     := '0';             --     peripheral_subsys_reset_in.reset_n
		sys_clk_timer_irq_irq                 : out std_logic                                         --              sys_clk_timer_irq.irq
	);
end entity peripheral_system;

architecture rtl of peripheral_system is
	component peripheral_system_button_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component peripheral_system_button_pio;

	component peripheral_system_high_res_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component peripheral_system_high_res_timer;

	component peripheral_system_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component peripheral_system_jtag_uart;

	component peripheral_system_led_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component peripheral_system_led_pio;

	component peripheral_system_performance_counter is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			write         : in  std_logic                     := 'X';             -- write
			writedata     : in  std_logic_vector(31 downto 0) := (others => 'X')  -- writedata
		);
	end component peripheral_system_performance_counter;

	component altera_avalon_mm_bridge is
		generic (
			DATA_WIDTH        : integer := 32;
			SYMBOL_WIDTH      : integer := 8;
			HDL_ADDR_WIDTH    : integer := 10;
			BURSTCOUNT_WIDTH  : integer := 1;
			PIPELINE_COMMAND  : integer := 1;
			PIPELINE_RESPONSE : integer := 1
		);
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset            : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(7 downto 0);                     -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic;                                        -- debugaccess
			s0_response      : out std_logic_vector(1 downto 0);                     -- response
			m0_response      : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- response
		);
	end component altera_avalon_mm_bridge;

	component peripheral_system_sys_clk_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component peripheral_system_sys_clk_timer;

	component peripheral_system_mm_interconnect_0 is
		port (
			clk_clk_clk                                         : in  std_logic                     := 'X';             -- clk
			peripheral_bridge_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			peripheral_bridge_m0_address                        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			peripheral_bridge_m0_waitrequest                    : out std_logic;                                        -- waitrequest
			peripheral_bridge_m0_burstcount                     : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			peripheral_bridge_m0_byteenable                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			peripheral_bridge_m0_read                           : in  std_logic                     := 'X';             -- read
			peripheral_bridge_m0_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			peripheral_bridge_m0_readdatavalid                  : out std_logic;                                        -- readdatavalid
			peripheral_bridge_m0_write                          : in  std_logic                     := 'X';             -- write
			peripheral_bridge_m0_writedata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			peripheral_bridge_m0_debugaccess                    : in  std_logic                     := 'X';             -- debugaccess
			button_pio_s1_address                               : out std_logic_vector(1 downto 0);                     -- address
			button_pio_s1_write                                 : out std_logic;                                        -- write
			button_pio_s1_readdata                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			button_pio_s1_writedata                             : out std_logic_vector(31 downto 0);                    -- writedata
			button_pio_s1_chipselect                            : out std_logic;                                        -- chipselect
			high_res_timer_s1_address                           : out std_logic_vector(2 downto 0);                     -- address
			high_res_timer_s1_write                             : out std_logic;                                        -- write
			high_res_timer_s1_readdata                          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			high_res_timer_s1_writedata                         : out std_logic_vector(15 downto 0);                    -- writedata
			high_res_timer_s1_chipselect                        : out std_logic;                                        -- chipselect
			jtag_uart_avalon_jtag_slave_address                 : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                   : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                    : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata               : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest             : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect              : out std_logic;                                        -- chipselect
			led_pio_s1_address                                  : out std_logic_vector(1 downto 0);                     -- address
			led_pio_s1_write                                    : out std_logic;                                        -- write
			led_pio_s1_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			led_pio_s1_writedata                                : out std_logic_vector(31 downto 0);                    -- writedata
			led_pio_s1_chipselect                               : out std_logic;                                        -- chipselect
			performance_counter_control_slave_address           : out std_logic_vector(3 downto 0);                     -- address
			performance_counter_control_slave_write             : out std_logic;                                        -- write
			performance_counter_control_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			performance_counter_control_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			performance_counter_control_slave_begintransfer     : out std_logic;                                        -- begintransfer
			sys_clk_timer_s1_address                            : out std_logic_vector(2 downto 0);                     -- address
			sys_clk_timer_s1_write                              : out std_logic;                                        -- write
			sys_clk_timer_s1_readdata                           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sys_clk_timer_s1_writedata                          : out std_logic_vector(15 downto 0);                    -- writedata
			sys_clk_timer_s1_chipselect                         : out std_logic                                         -- chipselect
		);
	end component peripheral_system_mm_interconnect_0;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal peripheral_bridge_m0_waitrequest                                  : std_logic;                     -- mm_interconnect_0:peripheral_bridge_m0_waitrequest -> peripheral_bridge:m0_waitrequest
	signal peripheral_bridge_m0_readdata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:peripheral_bridge_m0_readdata -> peripheral_bridge:m0_readdata
	signal peripheral_bridge_m0_debugaccess                                  : std_logic;                     -- peripheral_bridge:m0_debugaccess -> mm_interconnect_0:peripheral_bridge_m0_debugaccess
	signal peripheral_bridge_m0_address                                      : std_logic_vector(7 downto 0);  -- peripheral_bridge:m0_address -> mm_interconnect_0:peripheral_bridge_m0_address
	signal peripheral_bridge_m0_read                                         : std_logic;                     -- peripheral_bridge:m0_read -> mm_interconnect_0:peripheral_bridge_m0_read
	signal peripheral_bridge_m0_byteenable                                   : std_logic_vector(3 downto 0);  -- peripheral_bridge:m0_byteenable -> mm_interconnect_0:peripheral_bridge_m0_byteenable
	signal peripheral_bridge_m0_readdatavalid                                : std_logic;                     -- mm_interconnect_0:peripheral_bridge_m0_readdatavalid -> peripheral_bridge:m0_readdatavalid
	signal peripheral_bridge_m0_writedata                                    : std_logic_vector(31 downto 0); -- peripheral_bridge:m0_writedata -> mm_interconnect_0:peripheral_bridge_m0_writedata
	signal peripheral_bridge_m0_write                                        : std_logic;                     -- peripheral_bridge:m0_write -> mm_interconnect_0:peripheral_bridge_m0_write
	signal peripheral_bridge_m0_burstcount                                   : std_logic_vector(0 downto 0);  -- peripheral_bridge:m0_burstcount -> mm_interconnect_0:peripheral_bridge_m0_burstcount
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect          : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata            : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest         : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address             : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read                : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write               : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata           : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_performance_counter_control_slave_readdata      : std_logic_vector(31 downto 0); -- performance_counter:readdata -> mm_interconnect_0:performance_counter_control_slave_readdata
	signal mm_interconnect_0_performance_counter_control_slave_address       : std_logic_vector(3 downto 0);  -- mm_interconnect_0:performance_counter_control_slave_address -> performance_counter:address
	signal mm_interconnect_0_performance_counter_control_slave_begintransfer : std_logic;                     -- mm_interconnect_0:performance_counter_control_slave_begintransfer -> performance_counter:begintransfer
	signal mm_interconnect_0_performance_counter_control_slave_write         : std_logic;                     -- mm_interconnect_0:performance_counter_control_slave_write -> performance_counter:write
	signal mm_interconnect_0_performance_counter_control_slave_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:performance_counter_control_slave_writedata -> performance_counter:writedata
	signal mm_interconnect_0_sys_clk_timer_s1_chipselect                     : std_logic;                     -- mm_interconnect_0:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	signal mm_interconnect_0_sys_clk_timer_s1_readdata                       : std_logic_vector(15 downto 0); -- sys_clk_timer:readdata -> mm_interconnect_0:sys_clk_timer_s1_readdata
	signal mm_interconnect_0_sys_clk_timer_s1_address                        : std_logic_vector(2 downto 0);  -- mm_interconnect_0:sys_clk_timer_s1_address -> sys_clk_timer:address
	signal mm_interconnect_0_sys_clk_timer_s1_write                          : std_logic;                     -- mm_interconnect_0:sys_clk_timer_s1_write -> mm_interconnect_0_sys_clk_timer_s1_write:in
	signal mm_interconnect_0_sys_clk_timer_s1_writedata                      : std_logic_vector(15 downto 0); -- mm_interconnect_0:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	signal mm_interconnect_0_high_res_timer_s1_chipselect                    : std_logic;                     -- mm_interconnect_0:high_res_timer_s1_chipselect -> high_res_timer:chipselect
	signal mm_interconnect_0_high_res_timer_s1_readdata                      : std_logic_vector(15 downto 0); -- high_res_timer:readdata -> mm_interconnect_0:high_res_timer_s1_readdata
	signal mm_interconnect_0_high_res_timer_s1_address                       : std_logic_vector(2 downto 0);  -- mm_interconnect_0:high_res_timer_s1_address -> high_res_timer:address
	signal mm_interconnect_0_high_res_timer_s1_write                         : std_logic;                     -- mm_interconnect_0:high_res_timer_s1_write -> mm_interconnect_0_high_res_timer_s1_write:in
	signal mm_interconnect_0_high_res_timer_s1_writedata                     : std_logic_vector(15 downto 0); -- mm_interconnect_0:high_res_timer_s1_writedata -> high_res_timer:writedata
	signal mm_interconnect_0_button_pio_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:button_pio_s1_chipselect -> button_pio:chipselect
	signal mm_interconnect_0_button_pio_s1_readdata                          : std_logic_vector(31 downto 0); -- button_pio:readdata -> mm_interconnect_0:button_pio_s1_readdata
	signal mm_interconnect_0_button_pio_s1_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:button_pio_s1_address -> button_pio:address
	signal mm_interconnect_0_button_pio_s1_write                             : std_logic;                     -- mm_interconnect_0:button_pio_s1_write -> mm_interconnect_0_button_pio_s1_write:in
	signal mm_interconnect_0_button_pio_s1_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:button_pio_s1_writedata -> button_pio:writedata
	signal mm_interconnect_0_led_pio_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:led_pio_s1_chipselect -> led_pio:chipselect
	signal mm_interconnect_0_led_pio_s1_readdata                             : std_logic_vector(31 downto 0); -- led_pio:readdata -> mm_interconnect_0:led_pio_s1_readdata
	signal mm_interconnect_0_led_pio_s1_address                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:led_pio_s1_address -> led_pio:address
	signal mm_interconnect_0_led_pio_s1_write                                : std_logic;                     -- mm_interconnect_0:led_pio_s1_write -> mm_interconnect_0_led_pio_s1_write:in
	signal mm_interconnect_0_led_pio_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:led_pio_s1_writedata -> led_pio:writedata
	signal rst_controller_reset_out_reset                                    : std_logic;                     -- rst_controller:reset_out -> [mm_interconnect_0:peripheral_bridge_reset_reset_bridge_in_reset_reset, peripheral_bridge:reset, rst_controller_reset_out_reset:in]
	signal peripheral_subsys_reset_in_reset_n_ports_inv                      : std_logic;                     -- peripheral_subsys_reset_in_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv      : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv     : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_sys_clk_timer_s1_write_ports_inv                : std_logic;                     -- mm_interconnect_0_sys_clk_timer_s1_write:inv -> sys_clk_timer:write_n
	signal mm_interconnect_0_high_res_timer_s1_write_ports_inv               : std_logic;                     -- mm_interconnect_0_high_res_timer_s1_write:inv -> high_res_timer:write_n
	signal mm_interconnect_0_button_pio_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_0_button_pio_s1_write:inv -> button_pio:write_n
	signal mm_interconnect_0_led_pio_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_led_pio_s1_write:inv -> led_pio:write_n
	signal rst_controller_reset_out_reset_ports_inv                          : std_logic;                     -- rst_controller_reset_out_reset:inv -> [button_pio:reset_n, high_res_timer:reset_n, jtag_uart:rst_n, led_pio:reset_n, performance_counter:reset_n, sys_clk_timer:reset_n]

begin

	button_pio : component peripheral_system_button_pio
		port map (
			clk        => peripheral_subsys_clk_in_clk,                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,        --               reset.reset_n
			address    => mm_interconnect_0_button_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_button_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_button_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_button_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_button_pio_s1_readdata,        --                    .readdata
			in_port    => button_pio_external_connection_export,           -- external_connection.export
			irq        => button_pio_irq_irq                               --                 irq.irq
		);

	high_res_timer : component peripheral_system_high_res_timer
		port map (
			clk        => peripheral_subsys_clk_in_clk,                        --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,            -- reset.reset_n
			address    => mm_interconnect_0_high_res_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_high_res_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_high_res_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_high_res_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_high_res_timer_s1_write_ports_inv, --      .write_n
			irq        => high_res_timer_irq_irq                               --   irq.irq
		);

	jtag_uart : component peripheral_system_jtag_uart
		port map (
			clk            => peripheral_subsys_clk_in_clk,                                  --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => jtag_uart_irq_irq                                              --               irq.irq
		);

	led_pio : component peripheral_system_led_pio
		port map (
			clk        => peripheral_subsys_clk_in_clk,                 --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_led_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_led_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_led_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_led_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_led_pio_s1_readdata,        --                    .readdata
			out_port   => led_pio_external_connection_export            -- external_connection.export
		);

	performance_counter : component peripheral_system_performance_counter
		port map (
			clk           => peripheral_subsys_clk_in_clk,                                      --           clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                          --         reset.reset_n
			address       => mm_interconnect_0_performance_counter_control_slave_address,       -- control_slave.address
			begintransfer => mm_interconnect_0_performance_counter_control_slave_begintransfer, --              .begintransfer
			readdata      => mm_interconnect_0_performance_counter_control_slave_readdata,      --              .readdata
			write         => mm_interconnect_0_performance_counter_control_slave_write,         --              .write
			writedata     => mm_interconnect_0_performance_counter_control_slave_writedata      --              .writedata
		);

	peripheral_bridge : component altera_avalon_mm_bridge
		generic map (
			DATA_WIDTH        => 32,
			SYMBOL_WIDTH      => 8,
			HDL_ADDR_WIDTH    => 8,
			BURSTCOUNT_WIDTH  => 1,
			PIPELINE_COMMAND  => 1,
			PIPELINE_RESPONSE => 1
		)
		port map (
			clk              => peripheral_subsys_clk_in_clk,       --   clk.clk
			reset            => rst_controller_reset_out_reset,     -- reset.reset
			s0_waitrequest   => peripheral_bridge_s0_waitrequest,   --    s0.waitrequest
			s0_readdata      => peripheral_bridge_s0_readdata,      --      .readdata
			s0_readdatavalid => peripheral_bridge_s0_readdatavalid, --      .readdatavalid
			s0_burstcount    => peripheral_bridge_s0_burstcount,    --      .burstcount
			s0_writedata     => peripheral_bridge_s0_writedata,     --      .writedata
			s0_address       => peripheral_bridge_s0_address,       --      .address
			s0_write         => peripheral_bridge_s0_write,         --      .write
			s0_read          => peripheral_bridge_s0_read,          --      .read
			s0_byteenable    => peripheral_bridge_s0_byteenable,    --      .byteenable
			s0_debugaccess   => peripheral_bridge_s0_debugaccess,   --      .debugaccess
			m0_waitrequest   => peripheral_bridge_m0_waitrequest,   --    m0.waitrequest
			m0_readdata      => peripheral_bridge_m0_readdata,      --      .readdata
			m0_readdatavalid => peripheral_bridge_m0_readdatavalid, --      .readdatavalid
			m0_burstcount    => peripheral_bridge_m0_burstcount,    --      .burstcount
			m0_writedata     => peripheral_bridge_m0_writedata,     --      .writedata
			m0_address       => peripheral_bridge_m0_address,       --      .address
			m0_write         => peripheral_bridge_m0_write,         --      .write
			m0_read          => peripheral_bridge_m0_read,          --      .read
			m0_byteenable    => peripheral_bridge_m0_byteenable,    --      .byteenable
			m0_debugaccess   => peripheral_bridge_m0_debugaccess,   --      .debugaccess
			s0_response      => open,                               -- (terminated)
			m0_response      => "00"                                -- (terminated)
		);

	sys_clk_timer : component peripheral_system_sys_clk_timer
		port map (
			clk        => peripheral_subsys_clk_in_clk,                       --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,           -- reset.reset_n
			address    => mm_interconnect_0_sys_clk_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_sys_clk_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_sys_clk_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_sys_clk_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_sys_clk_timer_s1_write_ports_inv, --      .write_n
			irq        => sys_clk_timer_irq_irq                               --   irq.irq
		);

	mm_interconnect_0 : component peripheral_system_mm_interconnect_0
		port map (
			clk_clk_clk                                         => peripheral_subsys_clk_in_clk,                                      --                                       clk_clk.clk
			peripheral_bridge_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                                    -- peripheral_bridge_reset_reset_bridge_in_reset.reset
			peripheral_bridge_m0_address                        => peripheral_bridge_m0_address,                                      --                          peripheral_bridge_m0.address
			peripheral_bridge_m0_waitrequest                    => peripheral_bridge_m0_waitrequest,                                  --                                              .waitrequest
			peripheral_bridge_m0_burstcount                     => peripheral_bridge_m0_burstcount,                                   --                                              .burstcount
			peripheral_bridge_m0_byteenable                     => peripheral_bridge_m0_byteenable,                                   --                                              .byteenable
			peripheral_bridge_m0_read                           => peripheral_bridge_m0_read,                                         --                                              .read
			peripheral_bridge_m0_readdata                       => peripheral_bridge_m0_readdata,                                     --                                              .readdata
			peripheral_bridge_m0_readdatavalid                  => peripheral_bridge_m0_readdatavalid,                                --                                              .readdatavalid
			peripheral_bridge_m0_write                          => peripheral_bridge_m0_write,                                        --                                              .write
			peripheral_bridge_m0_writedata                      => peripheral_bridge_m0_writedata,                                    --                                              .writedata
			peripheral_bridge_m0_debugaccess                    => peripheral_bridge_m0_debugaccess,                                  --                                              .debugaccess
			button_pio_s1_address                               => mm_interconnect_0_button_pio_s1_address,                           --                                 button_pio_s1.address
			button_pio_s1_write                                 => mm_interconnect_0_button_pio_s1_write,                             --                                              .write
			button_pio_s1_readdata                              => mm_interconnect_0_button_pio_s1_readdata,                          --                                              .readdata
			button_pio_s1_writedata                             => mm_interconnect_0_button_pio_s1_writedata,                         --                                              .writedata
			button_pio_s1_chipselect                            => mm_interconnect_0_button_pio_s1_chipselect,                        --                                              .chipselect
			high_res_timer_s1_address                           => mm_interconnect_0_high_res_timer_s1_address,                       --                             high_res_timer_s1.address
			high_res_timer_s1_write                             => mm_interconnect_0_high_res_timer_s1_write,                         --                                              .write
			high_res_timer_s1_readdata                          => mm_interconnect_0_high_res_timer_s1_readdata,                      --                                              .readdata
			high_res_timer_s1_writedata                         => mm_interconnect_0_high_res_timer_s1_writedata,                     --                                              .writedata
			high_res_timer_s1_chipselect                        => mm_interconnect_0_high_res_timer_s1_chipselect,                    --                                              .chipselect
			jtag_uart_avalon_jtag_slave_address                 => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,             --                   jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,               --                                              .write
			jtag_uart_avalon_jtag_slave_read                    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,                --                                              .read
			jtag_uart_avalon_jtag_slave_readdata                => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,            --                                              .readdata
			jtag_uart_avalon_jtag_slave_writedata               => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,           --                                              .writedata
			jtag_uart_avalon_jtag_slave_waitrequest             => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,         --                                              .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect              => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,          --                                              .chipselect
			led_pio_s1_address                                  => mm_interconnect_0_led_pio_s1_address,                              --                                    led_pio_s1.address
			led_pio_s1_write                                    => mm_interconnect_0_led_pio_s1_write,                                --                                              .write
			led_pio_s1_readdata                                 => mm_interconnect_0_led_pio_s1_readdata,                             --                                              .readdata
			led_pio_s1_writedata                                => mm_interconnect_0_led_pio_s1_writedata,                            --                                              .writedata
			led_pio_s1_chipselect                               => mm_interconnect_0_led_pio_s1_chipselect,                           --                                              .chipselect
			performance_counter_control_slave_address           => mm_interconnect_0_performance_counter_control_slave_address,       --             performance_counter_control_slave.address
			performance_counter_control_slave_write             => mm_interconnect_0_performance_counter_control_slave_write,         --                                              .write
			performance_counter_control_slave_readdata          => mm_interconnect_0_performance_counter_control_slave_readdata,      --                                              .readdata
			performance_counter_control_slave_writedata         => mm_interconnect_0_performance_counter_control_slave_writedata,     --                                              .writedata
			performance_counter_control_slave_begintransfer     => mm_interconnect_0_performance_counter_control_slave_begintransfer, --                                              .begintransfer
			sys_clk_timer_s1_address                            => mm_interconnect_0_sys_clk_timer_s1_address,                        --                              sys_clk_timer_s1.address
			sys_clk_timer_s1_write                              => mm_interconnect_0_sys_clk_timer_s1_write,                          --                                              .write
			sys_clk_timer_s1_readdata                           => mm_interconnect_0_sys_clk_timer_s1_readdata,                       --                                              .readdata
			sys_clk_timer_s1_writedata                          => mm_interconnect_0_sys_clk_timer_s1_writedata,                      --                                              .writedata
			sys_clk_timer_s1_chipselect                         => mm_interconnect_0_sys_clk_timer_s1_chipselect                      --                                              .chipselect
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => peripheral_subsys_reset_in_reset_n_ports_inv, -- reset_in0.reset
			clk            => peripheral_subsys_clk_in_clk,                 --       clk.clk
			reset_out      => rst_controller_reset_out_reset,               -- reset_out.reset
			reset_req      => open,                                         -- (terminated)
			reset_req_in0  => '0',                                          -- (terminated)
			reset_in1      => '0',                                          -- (terminated)
			reset_req_in1  => '0',                                          -- (terminated)
			reset_in2      => '0',                                          -- (terminated)
			reset_req_in2  => '0',                                          -- (terminated)
			reset_in3      => '0',                                          -- (terminated)
			reset_req_in3  => '0',                                          -- (terminated)
			reset_in4      => '0',                                          -- (terminated)
			reset_req_in4  => '0',                                          -- (terminated)
			reset_in5      => '0',                                          -- (terminated)
			reset_req_in5  => '0',                                          -- (terminated)
			reset_in6      => '0',                                          -- (terminated)
			reset_req_in6  => '0',                                          -- (terminated)
			reset_in7      => '0',                                          -- (terminated)
			reset_req_in7  => '0',                                          -- (terminated)
			reset_in8      => '0',                                          -- (terminated)
			reset_req_in8  => '0',                                          -- (terminated)
			reset_in9      => '0',                                          -- (terminated)
			reset_req_in9  => '0',                                          -- (terminated)
			reset_in10     => '0',                                          -- (terminated)
			reset_req_in10 => '0',                                          -- (terminated)
			reset_in11     => '0',                                          -- (terminated)
			reset_req_in11 => '0',                                          -- (terminated)
			reset_in12     => '0',                                          -- (terminated)
			reset_req_in12 => '0',                                          -- (terminated)
			reset_in13     => '0',                                          -- (terminated)
			reset_req_in13 => '0',                                          -- (terminated)
			reset_in14     => '0',                                          -- (terminated)
			reset_req_in14 => '0',                                          -- (terminated)
			reset_in15     => '0',                                          -- (terminated)
			reset_req_in15 => '0'                                           -- (terminated)
		);

	peripheral_subsys_reset_in_reset_n_ports_inv <= not peripheral_subsys_reset_in_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_sys_clk_timer_s1_write_ports_inv <= not mm_interconnect_0_sys_clk_timer_s1_write;

	mm_interconnect_0_high_res_timer_s1_write_ports_inv <= not mm_interconnect_0_high_res_timer_s1_write;

	mm_interconnect_0_button_pio_s1_write_ports_inv <= not mm_interconnect_0_button_pio_s1_write;

	mm_interconnect_0_led_pio_s1_write_ports_inv <= not mm_interconnect_0_led_pio_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of peripheral_system
