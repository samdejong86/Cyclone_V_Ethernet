-- Nios_CPU_qsys.vhd

-- Generated using ACDS version 16.1 196

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Nios_CPU_qsys is
	port (
		clk_clk                                                    : in    std_logic                     := '0';             --                                 clk.clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_mem_clk               : out   std_logic;                                        --    mem_if_lpddr2_emif_0_pll_sharing.pll_mem_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_write_clk             : out   std_logic;                                        --                                    .pll_write_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_locked                : out   std_logic;                                        --                                    .pll_locked
		mem_if_lpddr2_emif_0_pll_sharing_pll_write_clk_pre_phy_clk : out   std_logic;                                        --                                    .pll_write_clk_pre_phy_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_addr_cmd_clk          : out   std_logic;                                        --                                    .pll_addr_cmd_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_avl_clk               : out   std_logic;                                        --                                    .pll_avl_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_config_clk            : out   std_logic;                                        --                                    .pll_config_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_mem_phy_clk           : out   std_logic;                                        --                                    .pll_mem_phy_clk
		mem_if_lpddr2_emif_0_pll_sharing_afi_phy_clk               : out   std_logic;                                        --                                    .afi_phy_clk
		mem_if_lpddr2_emif_0_pll_sharing_pll_avl_phy_clk           : out   std_logic;                                        --                                    .pll_avl_phy_clk
		mem_if_lpddr2_emif_0_status_local_init_done                : out   std_logic;                                        --         mem_if_lpddr2_emif_0_status.local_init_done
		mem_if_lpddr2_emif_0_status_local_cal_success              : out   std_logic;                                        --                                    .local_cal_success
		mem_if_lpddr2_emif_0_status_local_cal_fail                 : out   std_logic;                                        --                                    .local_cal_fail
		memory_mem_ca                                              : out   std_logic_vector(9 downto 0);                     --                              memory.mem_ca
		memory_mem_ck                                              : out   std_logic_vector(0 downto 0);                     --                                    .mem_ck
		memory_mem_ck_n                                            : out   std_logic_vector(0 downto 0);                     --                                    .mem_ck_n
		memory_mem_cke                                             : out   std_logic_vector(0 downto 0);                     --                                    .mem_cke
		memory_mem_cs_n                                            : out   std_logic_vector(0 downto 0);                     --                                    .mem_cs_n
		memory_mem_dm                                              : out   std_logic_vector(3 downto 0);                     --                                    .mem_dm
		memory_mem_dq                                              : inout std_logic_vector(31 downto 0) := (others => '0'); --                                    .mem_dq
		memory_mem_dqs                                             : inout std_logic_vector(3 downto 0)  := (others => '0'); --                                    .mem_dqs
		memory_mem_dqs_n                                           : inout std_logic_vector(3 downto 0)  := (others => '0'); --                                    .mem_dqs_n
		merged_resets_in_reset_reset_n                             : in    std_logic                     := '0';             --              merged_resets_in_reset.reset_n
		oct_rzqin                                                  : in    std_logic                     := '0';             --                                 oct.rzqin
		tse_mac_mac_gmii_connection_gmii_rx_d                      : in    std_logic_vector(7 downto 0)  := (others => '0'); --         tse_mac_mac_gmii_connection.gmii_rx_d
		tse_mac_mac_gmii_connection_gmii_rx_dv                     : in    std_logic                     := '0';             --                                    .gmii_rx_dv
		tse_mac_mac_gmii_connection_gmii_rx_err                    : in    std_logic                     := '0';             --                                    .gmii_rx_err
		tse_mac_mac_gmii_connection_gmii_tx_d                      : out   std_logic_vector(7 downto 0);                     --                                    .gmii_tx_d
		tse_mac_mac_gmii_connection_gmii_tx_en                     : out   std_logic;                                        --                                    .gmii_tx_en
		tse_mac_mac_gmii_connection_gmii_tx_err                    : out   std_logic;                                        --                                    .gmii_tx_err
		tse_mac_mac_mdio_connection_mdc                            : out   std_logic;                                        --         tse_mac_mac_mdio_connection.mdc
		tse_mac_mac_mdio_connection_mdio_in                        : in    std_logic                     := '0';             --                                    .mdio_in
		tse_mac_mac_mdio_connection_mdio_out                       : out   std_logic;                                        --                                    .mdio_out
		tse_mac_mac_mdio_connection_mdio_oen                       : out   std_logic;                                        --                                    .mdio_oen
		tse_mac_mac_mii_connection_mii_rx_d                        : in    std_logic_vector(3 downto 0)  := (others => '0'); --          tse_mac_mac_mii_connection.mii_rx_d
		tse_mac_mac_mii_connection_mii_rx_dv                       : in    std_logic                     := '0';             --                                    .mii_rx_dv
		tse_mac_mac_mii_connection_mii_rx_err                      : in    std_logic                     := '0';             --                                    .mii_rx_err
		tse_mac_mac_mii_connection_mii_tx_d                        : out   std_logic_vector(3 downto 0);                     --                                    .mii_tx_d
		tse_mac_mac_mii_connection_mii_tx_en                       : out   std_logic;                                        --                                    .mii_tx_en
		tse_mac_mac_mii_connection_mii_tx_err                      : out   std_logic;                                        --                                    .mii_tx_err
		tse_mac_mac_mii_connection_mii_crs                         : in    std_logic                     := '0';             --                                    .mii_crs
		tse_mac_mac_mii_connection_mii_col                         : in    std_logic                     := '0';             --                                    .mii_col
		tse_mac_mac_misc_connection_xon_gen                        : in    std_logic                     := '0';             --         tse_mac_mac_misc_connection.xon_gen
		tse_mac_mac_misc_connection_xoff_gen                       : in    std_logic                     := '0';             --                                    .xoff_gen
		tse_mac_mac_misc_connection_ff_tx_crc_fwd                  : in    std_logic                     := '0';             --                                    .ff_tx_crc_fwd
		tse_mac_mac_misc_connection_ff_tx_septy                    : out   std_logic;                                        --                                    .ff_tx_septy
		tse_mac_mac_misc_connection_tx_ff_uflow                    : out   std_logic;                                        --                                    .tx_ff_uflow
		tse_mac_mac_misc_connection_ff_tx_a_full                   : out   std_logic;                                        --                                    .ff_tx_a_full
		tse_mac_mac_misc_connection_ff_tx_a_empty                  : out   std_logic;                                        --                                    .ff_tx_a_empty
		tse_mac_mac_misc_connection_rx_err_stat                    : out   std_logic_vector(17 downto 0);                    --                                    .rx_err_stat
		tse_mac_mac_misc_connection_rx_frm_type                    : out   std_logic_vector(3 downto 0);                     --                                    .rx_frm_type
		tse_mac_mac_misc_connection_ff_rx_dsav                     : out   std_logic;                                        --                                    .ff_rx_dsav
		tse_mac_mac_misc_connection_ff_rx_a_full                   : out   std_logic;                                        --                                    .ff_rx_a_full
		tse_mac_mac_misc_connection_ff_rx_a_empty                  : out   std_logic;                                        --                                    .ff_rx_a_empty
		tse_mac_mac_status_connection_set_10                       : in    std_logic                     := '0';             --       tse_mac_mac_status_connection.set_10
		tse_mac_mac_status_connection_set_1000                     : in    std_logic                     := '0';             --                                    .set_1000
		tse_mac_mac_status_connection_eth_mode                     : out   std_logic;                                        --                                    .eth_mode
		tse_mac_mac_status_connection_ena_10                       : out   std_logic;                                        --                                    .ena_10
		tse_mac_pcs_mac_rx_clock_connection_clk                    : in    std_logic                     := '0';             -- tse_mac_pcs_mac_rx_clock_connection.clk
		tse_mac_pcs_mac_tx_clock_connection_clk                    : in    std_logic                     := '0'              -- tse_mac_pcs_mac_tx_clock_connection.clk
	);
end entity Nios_CPU_qsys;

architecture rtl of Nios_CPU_qsys is
	component Nios_CPU_qsys_cpu is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(30 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(30 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component Nios_CPU_qsys_cpu;

	component Nios_CPU_qsys_descriptor_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(10 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component Nios_CPU_qsys_descriptor_memory;

	component Nios_CPU_qsys_high_res_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component Nios_CPU_qsys_high_res_timer;

	component Nios_CPU_qsys_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component Nios_CPU_qsys_jtag_uart_0;

	component Nios_CPU_qsys_mem_if_lpddr2_emif_0 is
		port (
			pll_ref_clk                : in    std_logic                     := 'X';             -- clk
			global_reset_n             : in    std_logic                     := 'X';             -- reset_n
			soft_reset_n               : in    std_logic                     := 'X';             -- reset_n
			afi_clk                    : out   std_logic;                                        -- clk
			afi_half_clk               : out   std_logic;                                        -- clk
			afi_reset_n                : out   std_logic;                                        -- reset_n
			afi_reset_export_n         : out   std_logic;                                        -- reset_n
			mem_ca                     : out   std_logic_vector(9 downto 0);                     -- mem_ca
			mem_ck                     : out   std_logic_vector(0 downto 0);                     -- mem_ck
			mem_ck_n                   : out   std_logic_vector(0 downto 0);                     -- mem_ck_n
			mem_cke                    : out   std_logic_vector(0 downto 0);                     -- mem_cke
			mem_cs_n                   : out   std_logic_vector(0 downto 0);                     -- mem_cs_n
			mem_dm                     : out   std_logic_vector(3 downto 0);                     -- mem_dm
			mem_dq                     : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs                    : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n                  : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			avl_ready_0                : out   std_logic;                                        -- waitrequest_n
			avl_burstbegin_0           : in    std_logic                     := 'X';             -- beginbursttransfer
			avl_addr_0                 : in    std_logic_vector(26 downto 0) := (others => 'X'); -- address
			avl_rdata_valid_0          : out   std_logic;                                        -- readdatavalid
			avl_rdata_0                : out   std_logic_vector(31 downto 0);                    -- readdata
			avl_wdata_0                : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avl_be_0                   : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avl_read_req_0             : in    std_logic                     := 'X';             -- read
			avl_write_req_0            : in    std_logic                     := 'X';             -- write
			avl_size_0                 : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			mp_cmd_clk_0_clk           : in    std_logic                     := 'X';             -- clk
			mp_cmd_reset_n_0_reset_n   : in    std_logic                     := 'X';             -- reset_n
			mp_rfifo_clk_0_clk         : in    std_logic                     := 'X';             -- clk
			mp_rfifo_reset_n_0_reset_n : in    std_logic                     := 'X';             -- reset_n
			mp_wfifo_clk_0_clk         : in    std_logic                     := 'X';             -- clk
			mp_wfifo_reset_n_0_reset_n : in    std_logic                     := 'X';             -- reset_n
			local_init_done            : out   std_logic;                                        -- local_init_done
			local_cal_success          : out   std_logic;                                        -- local_cal_success
			local_cal_fail             : out   std_logic;                                        -- local_cal_fail
			oct_rzqin                  : in    std_logic                     := 'X';             -- rzqin
			pll_mem_clk                : out   std_logic;                                        -- pll_mem_clk
			pll_write_clk              : out   std_logic;                                        -- pll_write_clk
			pll_locked                 : out   std_logic;                                        -- pll_locked
			pll_write_clk_pre_phy_clk  : out   std_logic;                                        -- pll_write_clk_pre_phy_clk
			pll_addr_cmd_clk           : out   std_logic;                                        -- pll_addr_cmd_clk
			pll_avl_clk                : out   std_logic;                                        -- pll_avl_clk
			pll_config_clk             : out   std_logic;                                        -- pll_config_clk
			pll_mem_phy_clk            : out   std_logic;                                        -- pll_mem_phy_clk
			afi_phy_clk                : out   std_logic;                                        -- afi_phy_clk
			pll_avl_phy_clk            : out   std_logic                                         -- pll_avl_phy_clk
		);
	end component Nios_CPU_qsys_mem_if_lpddr2_emif_0;

	component Nios_CPU_qsys_onchip_ram is
		port (
			clk         : in  std_logic                     := 'X';             -- clk
			address     : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			clken       : in  std_logic                     := 'X';             -- clken
			chipselect  : in  std_logic                     := 'X';             -- chipselect
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset       : in  std_logic                     := 'X';             -- reset
			reset_req   : in  std_logic                     := 'X';             -- reset_req
			address2    : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			chipselect2 : in  std_logic                     := 'X';             -- chipselect
			clken2      : in  std_logic                     := 'X';             -- clken
			write2      : in  std_logic                     := 'X';             -- write
			readdata2   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata2  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable2 : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			clk2        : in  std_logic                     := 'X';             -- clk
			reset2      : in  std_logic                     := 'X';             -- reset
			reset_req2  : in  std_logic                     := 'X';             -- reset_req
			freeze      : in  std_logic                     := 'X'              -- freeze
		);
	end component Nios_CPU_qsys_onchip_ram;

	component altera_avalon_mm_bridge is
		generic (
			DATA_WIDTH        : integer := 32;
			SYMBOL_WIDTH      : integer := 8;
			HDL_ADDR_WIDTH    : integer := 10;
			BURSTCOUNT_WIDTH  : integer := 1;
			PIPELINE_COMMAND  : integer := 1;
			PIPELINE_RESPONSE : integer := 1
		);
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset            : in  std_logic                     := 'X';             -- reset
			s0_waitrequest   : out std_logic;                                        -- waitrequest
			s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			s0_readdatavalid : out std_logic;                                        -- readdatavalid
			s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			s0_address       : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			s0_write         : in  std_logic                     := 'X';             -- write
			s0_read          : in  std_logic                     := 'X';             -- read
			s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			m0_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			m0_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			m0_burstcount    : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			m0_address       : out std_logic_vector(9 downto 0);                     -- address
			m0_write         : out std_logic;                                        -- write
			m0_read          : out std_logic;                                        -- read
			m0_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess   : out std_logic;                                        -- debugaccess
			s0_response      : out std_logic_vector(1 downto 0);                     -- response
			m0_response      : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- response
		);
	end component altera_avalon_mm_bridge;

	component Nios_CPU_qsys_sgdma_rx is
		port (
			clk                           : in  std_logic                     := 'X';             -- clk
			system_reset_n                : in  std_logic                     := 'X';             -- reset_n
			csr_chipselect                : in  std_logic                     := 'X';             -- chipselect
			csr_address                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			csr_read                      : in  std_logic                     := 'X';             -- read
			csr_write                     : in  std_logic                     := 'X';             -- write
			csr_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			csr_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			descriptor_read_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			descriptor_read_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			descriptor_read_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			descriptor_read_address       : out std_logic_vector(31 downto 0);                    -- address
			descriptor_read_read          : out std_logic;                                        -- read
			descriptor_write_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			descriptor_write_address      : out std_logic_vector(31 downto 0);                    -- address
			descriptor_write_write        : out std_logic;                                        -- write
			descriptor_write_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			csr_irq                       : out std_logic;                                        -- irq
			in_startofpacket              : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket                : in  std_logic                     := 'X';             -- endofpacket
			in_data                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_valid                      : in  std_logic                     := 'X';             -- valid
			in_ready                      : out std_logic;                                        -- ready
			in_empty                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			in_error                      : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- error
			m_write_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			m_write_address               : out std_logic_vector(31 downto 0);                    -- address
			m_write_write                 : out std_logic;                                        -- write
			m_write_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			m_write_byteenable            : out std_logic_vector(3 downto 0)                      -- byteenable
		);
	end component Nios_CPU_qsys_sgdma_rx;

	component Nios_CPU_qsys_sgdma_tx is
		port (
			clk                           : in  std_logic                     := 'X';             -- clk
			system_reset_n                : in  std_logic                     := 'X';             -- reset_n
			csr_chipselect                : in  std_logic                     := 'X';             -- chipselect
			csr_address                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			csr_read                      : in  std_logic                     := 'X';             -- read
			csr_write                     : in  std_logic                     := 'X';             -- write
			csr_writedata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			csr_readdata                  : out std_logic_vector(31 downto 0);                    -- readdata
			descriptor_read_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			descriptor_read_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			descriptor_read_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			descriptor_read_address       : out std_logic_vector(31 downto 0);                    -- address
			descriptor_read_read          : out std_logic;                                        -- read
			descriptor_write_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			descriptor_write_address      : out std_logic_vector(31 downto 0);                    -- address
			descriptor_write_write        : out std_logic;                                        -- write
			descriptor_write_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			csr_irq                       : out std_logic;                                        -- irq
			m_read_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m_read_readdatavalid          : in  std_logic                     := 'X';             -- readdatavalid
			m_read_waitrequest            : in  std_logic                     := 'X';             -- waitrequest
			m_read_address                : out std_logic_vector(31 downto 0);                    -- address
			m_read_read                   : out std_logic;                                        -- read
			out_data                      : out std_logic_vector(31 downto 0);                    -- data
			out_valid                     : out std_logic;                                        -- valid
			out_ready                     : in  std_logic                     := 'X';             -- ready
			out_endofpacket               : out std_logic;                                        -- endofpacket
			out_startofpacket             : out std_logic;                                        -- startofpacket
			out_empty                     : out std_logic_vector(1 downto 0);                     -- empty
			out_error                     : out std_logic                                         -- error
		);
	end component Nios_CPU_qsys_sgdma_tx;

	component Nios_CPU_qsys_sys_clk_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component Nios_CPU_qsys_sys_clk_timer;

	component Nios_CPU_qsys_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component Nios_CPU_qsys_sysid;

	component Nios_CPU_qsys_tse_mac is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			reg_addr      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			reg_data_out  : out std_logic_vector(31 downto 0);                    -- readdata
			reg_rd        : in  std_logic                     := 'X';             -- read
			reg_data_in   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			reg_wr        : in  std_logic                     := 'X';             -- write
			reg_busy      : out std_logic;                                        -- waitrequest
			tx_clk        : in  std_logic                     := 'X';             -- clk
			rx_clk        : in  std_logic                     := 'X';             -- clk
			set_10        : in  std_logic                     := 'X';             -- set_10
			set_1000      : in  std_logic                     := 'X';             -- set_1000
			eth_mode      : out std_logic;                                        -- eth_mode
			ena_10        : out std_logic;                                        -- ena_10
			gm_rx_d       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- gmii_rx_d
			gm_rx_dv      : in  std_logic                     := 'X';             -- gmii_rx_dv
			gm_rx_err     : in  std_logic                     := 'X';             -- gmii_rx_err
			gm_tx_d       : out std_logic_vector(7 downto 0);                     -- gmii_tx_d
			gm_tx_en      : out std_logic;                                        -- gmii_tx_en
			gm_tx_err     : out std_logic;                                        -- gmii_tx_err
			m_rx_d        : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- mii_rx_d
			m_rx_en       : in  std_logic                     := 'X';             -- mii_rx_dv
			m_rx_err      : in  std_logic                     := 'X';             -- mii_rx_err
			m_tx_d        : out std_logic_vector(3 downto 0);                     -- mii_tx_d
			m_tx_en       : out std_logic;                                        -- mii_tx_en
			m_tx_err      : out std_logic;                                        -- mii_tx_err
			m_rx_crs      : in  std_logic                     := 'X';             -- mii_crs
			m_rx_col      : in  std_logic                     := 'X';             -- mii_col
			ff_rx_clk     : in  std_logic                     := 'X';             -- clk
			ff_tx_clk     : in  std_logic                     := 'X';             -- clk
			ff_rx_data    : out std_logic_vector(31 downto 0);                    -- data
			ff_rx_eop     : out std_logic;                                        -- endofpacket
			rx_err        : out std_logic_vector(5 downto 0);                     -- error
			ff_rx_mod     : out std_logic_vector(1 downto 0);                     -- empty
			ff_rx_rdy     : in  std_logic                     := 'X';             -- ready
			ff_rx_sop     : out std_logic;                                        -- startofpacket
			ff_rx_dval    : out std_logic;                                        -- valid
			ff_tx_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			ff_tx_eop     : in  std_logic                     := 'X';             -- endofpacket
			ff_tx_err     : in  std_logic                     := 'X';             -- error
			ff_tx_mod     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			ff_tx_rdy     : out std_logic;                                        -- ready
			ff_tx_sop     : in  std_logic                     := 'X';             -- startofpacket
			ff_tx_wren    : in  std_logic                     := 'X';             -- valid
			mdc           : out std_logic;                                        -- mdc
			mdio_in       : in  std_logic                     := 'X';             -- mdio_in
			mdio_out      : out std_logic;                                        -- mdio_out
			mdio_oen      : out std_logic;                                        -- mdio_oen
			xon_gen       : in  std_logic                     := 'X';             -- xon_gen
			xoff_gen      : in  std_logic                     := 'X';             -- xoff_gen
			ff_tx_crc_fwd : in  std_logic                     := 'X';             -- ff_tx_crc_fwd
			ff_tx_septy   : out std_logic;                                        -- ff_tx_septy
			tx_ff_uflow   : out std_logic;                                        -- tx_ff_uflow
			ff_tx_a_full  : out std_logic;                                        -- ff_tx_a_full
			ff_tx_a_empty : out std_logic;                                        -- ff_tx_a_empty
			rx_err_stat   : out std_logic_vector(17 downto 0);                    -- rx_err_stat
			rx_frm_type   : out std_logic_vector(3 downto 0);                     -- rx_frm_type
			ff_rx_dsav    : out std_logic;                                        -- ff_rx_dsav
			ff_rx_a_full  : out std_logic;                                        -- ff_rx_a_full
			ff_rx_a_empty : out std_logic                                         -- ff_rx_a_empty
		);
	end component Nios_CPU_qsys_tse_mac;

	component Nios_CPU_qsys_mm_interconnect_0 is
		port (
			clkin_50_clk_clk                                                        : in  std_logic                     := 'X';             -- clk
			mem_if_lpddr2_emif_0_afi_clk_clk                                        : in  std_logic                     := 'X';             -- clk
			cpu_reset_reset_bridge_in_reset_reset                                   : in  std_logic                     := 'X';             -- reset
			mem_if_lpddr2_emif_0_avl_0_translator_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			mem_if_lpddr2_emif_0_mp_cmd_reset_n_0_reset_bridge_in_reset_reset       : in  std_logic                     := 'X';             -- reset
			sgdma_rx_reset_reset_bridge_in_reset_reset                              : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                                                 : in  std_logic_vector(30 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest                                             : out std_logic;                                        -- waitrequest
			cpu_data_master_byteenable                                              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                                                    : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                                                : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_readdatavalid                                           : out std_logic;                                        -- readdatavalid
			cpu_data_master_write                                                   : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata                                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess                                             : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address                                          : in  std_logic_vector(30 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest                                      : out std_logic;                                        -- waitrequest
			cpu_instruction_master_read                                             : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata                                         : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_instruction_master_readdatavalid                                    : out std_logic;                                        -- readdatavalid
			sgdma_rx_descriptor_read_address                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_rx_descriptor_read_waitrequest                                    : out std_logic;                                        -- waitrequest
			sgdma_rx_descriptor_read_read                                           : in  std_logic                     := 'X';             -- read
			sgdma_rx_descriptor_read_readdata                                       : out std_logic_vector(31 downto 0);                    -- readdata
			sgdma_rx_descriptor_read_readdatavalid                                  : out std_logic;                                        -- readdatavalid
			sgdma_rx_descriptor_write_address                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_rx_descriptor_write_waitrequest                                   : out std_logic;                                        -- waitrequest
			sgdma_rx_descriptor_write_write                                         : in  std_logic                     := 'X';             -- write
			sgdma_rx_descriptor_write_writedata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			sgdma_rx_m_write_address                                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_rx_m_write_waitrequest                                            : out std_logic;                                        -- waitrequest
			sgdma_rx_m_write_byteenable                                             : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			sgdma_rx_m_write_write                                                  : in  std_logic                     := 'X';             -- write
			sgdma_rx_m_write_writedata                                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			sgdma_tx_descriptor_read_address                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_tx_descriptor_read_waitrequest                                    : out std_logic;                                        -- waitrequest
			sgdma_tx_descriptor_read_read                                           : in  std_logic                     := 'X';             -- read
			sgdma_tx_descriptor_read_readdata                                       : out std_logic_vector(31 downto 0);                    -- readdata
			sgdma_tx_descriptor_read_readdatavalid                                  : out std_logic;                                        -- readdatavalid
			sgdma_tx_descriptor_write_address                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_tx_descriptor_write_waitrequest                                   : out std_logic;                                        -- waitrequest
			sgdma_tx_descriptor_write_write                                         : in  std_logic                     := 'X';             -- write
			sgdma_tx_descriptor_write_writedata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			sgdma_tx_m_read_address                                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			sgdma_tx_m_read_waitrequest                                             : out std_logic;                                        -- waitrequest
			sgdma_tx_m_read_read                                                    : in  std_logic                     := 'X';             -- read
			sgdma_tx_m_read_readdata                                                : out std_logic_vector(31 downto 0);                    -- readdata
			sgdma_tx_m_read_readdatavalid                                           : out std_logic;                                        -- readdatavalid
			cpu_debug_mem_slave_address                                             : out std_logic_vector(8 downto 0);                     -- address
			cpu_debug_mem_slave_write                                               : out std_logic;                                        -- write
			cpu_debug_mem_slave_read                                                : out std_logic;                                        -- read
			cpu_debug_mem_slave_readdata                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_debug_mem_slave_writedata                                           : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_debug_mem_slave_byteenable                                          : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_debug_mem_slave_waitrequest                                         : in  std_logic                     := 'X';             -- waitrequest
			cpu_debug_mem_slave_debugaccess                                         : out std_logic;                                        -- debugaccess
			descriptor_memory_s1_address                                            : out std_logic_vector(10 downto 0);                    -- address
			descriptor_memory_s1_write                                              : out std_logic;                                        -- write
			descriptor_memory_s1_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			descriptor_memory_s1_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			descriptor_memory_s1_byteenable                                         : out std_logic_vector(3 downto 0);                     -- byteenable
			descriptor_memory_s1_chipselect                                         : out std_logic;                                        -- chipselect
			descriptor_memory_s1_clken                                              : out std_logic;                                        -- clken
			mem_if_lpddr2_emif_0_avl_0_address                                      : out std_logic_vector(26 downto 0);                    -- address
			mem_if_lpddr2_emif_0_avl_0_write                                        : out std_logic;                                        -- write
			mem_if_lpddr2_emif_0_avl_0_read                                         : out std_logic;                                        -- read
			mem_if_lpddr2_emif_0_avl_0_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			mem_if_lpddr2_emif_0_avl_0_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			mem_if_lpddr2_emif_0_avl_0_beginbursttransfer                           : out std_logic;                                        -- beginbursttransfer
			mem_if_lpddr2_emif_0_avl_0_burstcount                                   : out std_logic_vector(2 downto 0);                     -- burstcount
			mem_if_lpddr2_emif_0_avl_0_byteenable                                   : out std_logic_vector(3 downto 0);                     -- byteenable
			mem_if_lpddr2_emif_0_avl_0_readdatavalid                                : in  std_logic                     := 'X';             -- readdatavalid
			mem_if_lpddr2_emif_0_avl_0_waitrequest                                  : in  std_logic                     := 'X';             -- waitrequest
			onchip_ram_s1_address                                                   : out std_logic_vector(18 downto 0);                    -- address
			onchip_ram_s1_write                                                     : out std_logic;                                        -- write
			onchip_ram_s1_readdata                                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_ram_s1_writedata                                                 : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_ram_s1_byteenable                                                : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_ram_s1_chipselect                                                : out std_logic;                                        -- chipselect
			onchip_ram_s1_clken                                                     : out std_logic;                                        -- clken
			onchip_ram_s2_address                                                   : out std_logic_vector(18 downto 0);                    -- address
			onchip_ram_s2_write                                                     : out std_logic;                                        -- write
			onchip_ram_s2_readdata                                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_ram_s2_writedata                                                 : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_ram_s2_byteenable                                                : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_ram_s2_chipselect                                                : out std_logic;                                        -- chipselect
			onchip_ram_s2_clken                                                     : out std_logic;                                        -- clken
			pb_cpu_to_io_s0_address                                                 : out std_logic_vector(9 downto 0);                     -- address
			pb_cpu_to_io_s0_write                                                   : out std_logic;                                        -- write
			pb_cpu_to_io_s0_read                                                    : out std_logic;                                        -- read
			pb_cpu_to_io_s0_readdata                                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pb_cpu_to_io_s0_writedata                                               : out std_logic_vector(31 downto 0);                    -- writedata
			pb_cpu_to_io_s0_burstcount                                              : out std_logic_vector(0 downto 0);                     -- burstcount
			pb_cpu_to_io_s0_byteenable                                              : out std_logic_vector(3 downto 0);                     -- byteenable
			pb_cpu_to_io_s0_readdatavalid                                           : in  std_logic                     := 'X';             -- readdatavalid
			pb_cpu_to_io_s0_waitrequest                                             : in  std_logic                     := 'X';             -- waitrequest
			pb_cpu_to_io_s0_debugaccess                                             : out std_logic;                                        -- debugaccess
			sgdma_rx_csr_address                                                    : out std_logic_vector(3 downto 0);                     -- address
			sgdma_rx_csr_write                                                      : out std_logic;                                        -- write
			sgdma_rx_csr_read                                                       : out std_logic;                                        -- read
			sgdma_rx_csr_readdata                                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sgdma_rx_csr_writedata                                                  : out std_logic_vector(31 downto 0);                    -- writedata
			sgdma_rx_csr_chipselect                                                 : out std_logic;                                        -- chipselect
			sgdma_tx_csr_address                                                    : out std_logic_vector(3 downto 0);                     -- address
			sgdma_tx_csr_write                                                      : out std_logic;                                        -- write
			sgdma_tx_csr_read                                                       : out std_logic;                                        -- read
			sgdma_tx_csr_readdata                                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sgdma_tx_csr_writedata                                                  : out std_logic_vector(31 downto 0);                    -- writedata
			sgdma_tx_csr_chipselect                                                 : out std_logic;                                        -- chipselect
			tse_mac_control_port_address                                            : out std_logic_vector(7 downto 0);                     -- address
			tse_mac_control_port_write                                              : out std_logic;                                        -- write
			tse_mac_control_port_read                                               : out std_logic;                                        -- read
			tse_mac_control_port_readdata                                           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			tse_mac_control_port_writedata                                          : out std_logic_vector(31 downto 0);                    -- writedata
			tse_mac_control_port_waitrequest                                        : in  std_logic                     := 'X'              -- waitrequest
		);
	end component Nios_CPU_qsys_mm_interconnect_0;

	component Nios_CPU_qsys_mm_interconnect_1 is
		port (
			clkin_50_clk_clk                               : in  std_logic                     := 'X';             -- clk
			jtag_uart_0_reset_reset_bridge_in_reset_reset  : in  std_logic                     := 'X';             -- reset
			pb_cpu_to_io_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			pb_cpu_to_io_m0_address                        : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			pb_cpu_to_io_m0_waitrequest                    : out std_logic;                                        -- waitrequest
			pb_cpu_to_io_m0_burstcount                     : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			pb_cpu_to_io_m0_byteenable                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			pb_cpu_to_io_m0_read                           : in  std_logic                     := 'X';             -- read
			pb_cpu_to_io_m0_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			pb_cpu_to_io_m0_readdatavalid                  : out std_logic;                                        -- readdatavalid
			pb_cpu_to_io_m0_write                          : in  std_logic                     := 'X';             -- write
			pb_cpu_to_io_m0_writedata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			pb_cpu_to_io_m0_debugaccess                    : in  std_logic                     := 'X';             -- debugaccess
			high_res_timer_s1_address                      : out std_logic_vector(2 downto 0);                     -- address
			high_res_timer_s1_write                        : out std_logic;                                        -- write
			high_res_timer_s1_readdata                     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			high_res_timer_s1_writedata                    : out std_logic_vector(15 downto 0);                    -- writedata
			high_res_timer_s1_chipselect                   : out std_logic;                                        -- chipselect
			jtag_uart_0_avalon_jtag_slave_address          : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write            : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read             : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest      : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect       : out std_logic;                                        -- chipselect
			sys_clk_timer_s1_address                       : out std_logic_vector(2 downto 0);                     -- address
			sys_clk_timer_s1_write                         : out std_logic;                                        -- write
			sys_clk_timer_s1_readdata                      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sys_clk_timer_s1_writedata                     : out std_logic_vector(15 downto 0);                    -- writedata
			sys_clk_timer_s1_chipselect                    : out std_logic;                                        -- chipselect
			sysid_control_slave_address                    : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component Nios_CPU_qsys_mm_interconnect_1;

	component Nios_CPU_qsys_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component Nios_CPU_qsys_irq_mapper;

	component Nios_CPU_qsys_avalon_st_adapter is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk        : in  std_logic                     := 'X';             -- clk
			in_rst_0_reset      : in  std_logic                     := 'X';             -- reset
			in_0_data           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			in_0_valid          : in  std_logic                     := 'X';             -- valid
			in_0_ready          : out std_logic;                                        -- ready
			in_0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			in_0_empty          : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- empty
			in_0_error          : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- error
			out_0_data          : out std_logic_vector(31 downto 0);                    -- data
			out_0_valid         : out std_logic;                                        -- valid
			out_0_ready         : in  std_logic                     := 'X';             -- ready
			out_0_startofpacket : out std_logic;                                        -- startofpacket
			out_0_endofpacket   : out std_logic;                                        -- endofpacket
			out_0_empty         : out std_logic_vector(1 downto 0);                     -- empty
			out_0_error         : out std_logic_vector(5 downto 0)                      -- error
		);
	end component Nios_CPU_qsys_avalon_st_adapter;

	component nios_cpu_qsys_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_in2      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component nios_cpu_qsys_rst_controller;

	component nios_cpu_qsys_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component nios_cpu_qsys_rst_controller_001;

	component nios_cpu_qsys_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component nios_cpu_qsys_rst_controller_002;

	signal sgdma_tx_out_valid                                              : std_logic;                     -- sgdma_tx:out_valid -> tse_mac:ff_tx_wren
	signal sgdma_tx_out_data                                               : std_logic_vector(31 downto 0); -- sgdma_tx:out_data -> tse_mac:ff_tx_data
	signal sgdma_tx_out_ready                                              : std_logic;                     -- tse_mac:ff_tx_rdy -> sgdma_tx:out_ready
	signal sgdma_tx_out_startofpacket                                      : std_logic;                     -- sgdma_tx:out_startofpacket -> tse_mac:ff_tx_sop
	signal sgdma_tx_out_endofpacket                                        : std_logic;                     -- sgdma_tx:out_endofpacket -> tse_mac:ff_tx_eop
	signal sgdma_tx_out_error                                              : std_logic;                     -- sgdma_tx:out_error -> tse_mac:ff_tx_err
	signal sgdma_tx_out_empty                                              : std_logic_vector(1 downto 0);  -- sgdma_tx:out_empty -> tse_mac:ff_tx_mod
	signal mem_if_lpddr2_emif_0_afi_clk_clk                                : std_logic;                     -- mem_if_lpddr2_emif_0:afi_clk -> [mem_if_lpddr2_emif_0:mp_cmd_clk_0_clk, mem_if_lpddr2_emif_0:mp_rfifo_clk_0_clk, mem_if_lpddr2_emif_0:mp_wfifo_clk_0_clk, mm_interconnect_0:mem_if_lpddr2_emif_0_afi_clk_clk, rst_controller_002:clk]
	signal cpu_data_master_readdata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_waitrequest                                     : std_logic;                     -- mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_debugaccess                                     : std_logic;                     -- cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	signal cpu_data_master_address                                         : std_logic_vector(30 downto 0); -- cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	signal cpu_data_master_byteenable                                      : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	signal cpu_data_master_read                                            : std_logic;                     -- cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	signal cpu_data_master_readdatavalid                                   : std_logic;                     -- mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	signal cpu_data_master_write                                           : std_logic;                     -- cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	signal cpu_data_master_writedata                                       : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	signal sgdma_rx_descriptor_read_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:sgdma_rx_descriptor_read_readdata -> sgdma_rx:descriptor_read_readdata
	signal sgdma_rx_descriptor_read_waitrequest                            : std_logic;                     -- mm_interconnect_0:sgdma_rx_descriptor_read_waitrequest -> sgdma_rx:descriptor_read_waitrequest
	signal sgdma_rx_descriptor_read_address                                : std_logic_vector(31 downto 0); -- sgdma_rx:descriptor_read_address -> mm_interconnect_0:sgdma_rx_descriptor_read_address
	signal sgdma_rx_descriptor_read_read                                   : std_logic;                     -- sgdma_rx:descriptor_read_read -> mm_interconnect_0:sgdma_rx_descriptor_read_read
	signal sgdma_rx_descriptor_read_readdatavalid                          : std_logic;                     -- mm_interconnect_0:sgdma_rx_descriptor_read_readdatavalid -> sgdma_rx:descriptor_read_readdatavalid
	signal cpu_instruction_master_readdata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_waitrequest                              : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                  : std_logic_vector(30 downto 0); -- cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	signal cpu_instruction_master_read                                     : std_logic;                     -- cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	signal cpu_instruction_master_readdatavalid                            : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	signal sgdma_tx_m_read_readdata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:sgdma_tx_m_read_readdata -> sgdma_tx:m_read_readdata
	signal sgdma_tx_m_read_waitrequest                                     : std_logic;                     -- mm_interconnect_0:sgdma_tx_m_read_waitrequest -> sgdma_tx:m_read_waitrequest
	signal sgdma_tx_m_read_address                                         : std_logic_vector(31 downto 0); -- sgdma_tx:m_read_address -> mm_interconnect_0:sgdma_tx_m_read_address
	signal sgdma_tx_m_read_read                                            : std_logic;                     -- sgdma_tx:m_read_read -> mm_interconnect_0:sgdma_tx_m_read_read
	signal sgdma_tx_m_read_readdatavalid                                   : std_logic;                     -- mm_interconnect_0:sgdma_tx_m_read_readdatavalid -> sgdma_tx:m_read_readdatavalid
	signal sgdma_rx_m_write_waitrequest                                    : std_logic;                     -- mm_interconnect_0:sgdma_rx_m_write_waitrequest -> sgdma_rx:m_write_waitrequest
	signal sgdma_rx_m_write_address                                        : std_logic_vector(31 downto 0); -- sgdma_rx:m_write_address -> mm_interconnect_0:sgdma_rx_m_write_address
	signal sgdma_rx_m_write_byteenable                                     : std_logic_vector(3 downto 0);  -- sgdma_rx:m_write_byteenable -> mm_interconnect_0:sgdma_rx_m_write_byteenable
	signal sgdma_rx_m_write_write                                          : std_logic;                     -- sgdma_rx:m_write_write -> mm_interconnect_0:sgdma_rx_m_write_write
	signal sgdma_rx_m_write_writedata                                      : std_logic_vector(31 downto 0); -- sgdma_rx:m_write_writedata -> mm_interconnect_0:sgdma_rx_m_write_writedata
	signal sgdma_tx_descriptor_read_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:sgdma_tx_descriptor_read_readdata -> sgdma_tx:descriptor_read_readdata
	signal sgdma_tx_descriptor_read_waitrequest                            : std_logic;                     -- mm_interconnect_0:sgdma_tx_descriptor_read_waitrequest -> sgdma_tx:descriptor_read_waitrequest
	signal sgdma_tx_descriptor_read_address                                : std_logic_vector(31 downto 0); -- sgdma_tx:descriptor_read_address -> mm_interconnect_0:sgdma_tx_descriptor_read_address
	signal sgdma_tx_descriptor_read_read                                   : std_logic;                     -- sgdma_tx:descriptor_read_read -> mm_interconnect_0:sgdma_tx_descriptor_read_read
	signal sgdma_tx_descriptor_read_readdatavalid                          : std_logic;                     -- mm_interconnect_0:sgdma_tx_descriptor_read_readdatavalid -> sgdma_tx:descriptor_read_readdatavalid
	signal sgdma_rx_descriptor_write_waitrequest                           : std_logic;                     -- mm_interconnect_0:sgdma_rx_descriptor_write_waitrequest -> sgdma_rx:descriptor_write_waitrequest
	signal sgdma_rx_descriptor_write_address                               : std_logic_vector(31 downto 0); -- sgdma_rx:descriptor_write_address -> mm_interconnect_0:sgdma_rx_descriptor_write_address
	signal sgdma_rx_descriptor_write_write                                 : std_logic;                     -- sgdma_rx:descriptor_write_write -> mm_interconnect_0:sgdma_rx_descriptor_write_write
	signal sgdma_rx_descriptor_write_writedata                             : std_logic_vector(31 downto 0); -- sgdma_rx:descriptor_write_writedata -> mm_interconnect_0:sgdma_rx_descriptor_write_writedata
	signal sgdma_tx_descriptor_write_waitrequest                           : std_logic;                     -- mm_interconnect_0:sgdma_tx_descriptor_write_waitrequest -> sgdma_tx:descriptor_write_waitrequest
	signal sgdma_tx_descriptor_write_address                               : std_logic_vector(31 downto 0); -- sgdma_tx:descriptor_write_address -> mm_interconnect_0:sgdma_tx_descriptor_write_address
	signal sgdma_tx_descriptor_write_write                                 : std_logic;                     -- sgdma_tx:descriptor_write_write -> mm_interconnect_0:sgdma_tx_descriptor_write_write
	signal sgdma_tx_descriptor_write_writedata                             : std_logic_vector(31 downto 0); -- sgdma_tx:descriptor_write_writedata -> mm_interconnect_0:sgdma_tx_descriptor_write_writedata
	signal mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_beginbursttransfer : std_logic;                     -- mm_interconnect_0:mem_if_lpddr2_emif_0_avl_0_beginbursttransfer -> mem_if_lpddr2_emif_0:avl_burstbegin_0
	signal mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_readdata           : std_logic_vector(31 downto 0); -- mem_if_lpddr2_emif_0:avl_rdata_0 -> mm_interconnect_0:mem_if_lpddr2_emif_0_avl_0_readdata
	signal mem_if_lpddr2_emif_0_avl_0_waitrequest                          : std_logic;                     -- mem_if_lpddr2_emif_0:avl_ready_0 -> mem_if_lpddr2_emif_0_avl_0_waitrequest:in
	signal mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_address            : std_logic_vector(26 downto 0); -- mm_interconnect_0:mem_if_lpddr2_emif_0_avl_0_address -> mem_if_lpddr2_emif_0:avl_addr_0
	signal mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_read               : std_logic;                     -- mm_interconnect_0:mem_if_lpddr2_emif_0_avl_0_read -> mem_if_lpddr2_emif_0:avl_read_req_0
	signal mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_byteenable         : std_logic_vector(3 downto 0);  -- mm_interconnect_0:mem_if_lpddr2_emif_0_avl_0_byteenable -> mem_if_lpddr2_emif_0:avl_be_0
	signal mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_readdatavalid      : std_logic;                     -- mem_if_lpddr2_emif_0:avl_rdata_valid_0 -> mm_interconnect_0:mem_if_lpddr2_emif_0_avl_0_readdatavalid
	signal mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_write              : std_logic;                     -- mm_interconnect_0:mem_if_lpddr2_emif_0_avl_0_write -> mem_if_lpddr2_emif_0:avl_write_req_0
	signal mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_writedata          : std_logic_vector(31 downto 0); -- mm_interconnect_0:mem_if_lpddr2_emif_0_avl_0_writedata -> mem_if_lpddr2_emif_0:avl_wdata_0
	signal mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_burstcount         : std_logic_vector(2 downto 0);  -- mm_interconnect_0:mem_if_lpddr2_emif_0_avl_0_burstcount -> mem_if_lpddr2_emif_0:avl_size_0
	signal mm_interconnect_0_tse_mac_control_port_readdata                 : std_logic_vector(31 downto 0); -- tse_mac:reg_data_out -> mm_interconnect_0:tse_mac_control_port_readdata
	signal mm_interconnect_0_tse_mac_control_port_waitrequest              : std_logic;                     -- tse_mac:reg_busy -> mm_interconnect_0:tse_mac_control_port_waitrequest
	signal mm_interconnect_0_tse_mac_control_port_address                  : std_logic_vector(7 downto 0);  -- mm_interconnect_0:tse_mac_control_port_address -> tse_mac:reg_addr
	signal mm_interconnect_0_tse_mac_control_port_read                     : std_logic;                     -- mm_interconnect_0:tse_mac_control_port_read -> tse_mac:reg_rd
	signal mm_interconnect_0_tse_mac_control_port_write                    : std_logic;                     -- mm_interconnect_0:tse_mac_control_port_write -> tse_mac:reg_wr
	signal mm_interconnect_0_tse_mac_control_port_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:tse_mac_control_port_writedata -> tse_mac:reg_data_in
	signal mm_interconnect_0_sgdma_tx_csr_chipselect                       : std_logic;                     -- mm_interconnect_0:sgdma_tx_csr_chipselect -> sgdma_tx:csr_chipselect
	signal mm_interconnect_0_sgdma_tx_csr_readdata                         : std_logic_vector(31 downto 0); -- sgdma_tx:csr_readdata -> mm_interconnect_0:sgdma_tx_csr_readdata
	signal mm_interconnect_0_sgdma_tx_csr_address                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:sgdma_tx_csr_address -> sgdma_tx:csr_address
	signal mm_interconnect_0_sgdma_tx_csr_read                             : std_logic;                     -- mm_interconnect_0:sgdma_tx_csr_read -> sgdma_tx:csr_read
	signal mm_interconnect_0_sgdma_tx_csr_write                            : std_logic;                     -- mm_interconnect_0:sgdma_tx_csr_write -> sgdma_tx:csr_write
	signal mm_interconnect_0_sgdma_tx_csr_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:sgdma_tx_csr_writedata -> sgdma_tx:csr_writedata
	signal mm_interconnect_0_sgdma_rx_csr_chipselect                       : std_logic;                     -- mm_interconnect_0:sgdma_rx_csr_chipselect -> sgdma_rx:csr_chipselect
	signal mm_interconnect_0_sgdma_rx_csr_readdata                         : std_logic_vector(31 downto 0); -- sgdma_rx:csr_readdata -> mm_interconnect_0:sgdma_rx_csr_readdata
	signal mm_interconnect_0_sgdma_rx_csr_address                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:sgdma_rx_csr_address -> sgdma_rx:csr_address
	signal mm_interconnect_0_sgdma_rx_csr_read                             : std_logic;                     -- mm_interconnect_0:sgdma_rx_csr_read -> sgdma_rx:csr_read
	signal mm_interconnect_0_sgdma_rx_csr_write                            : std_logic;                     -- mm_interconnect_0:sgdma_rx_csr_write -> sgdma_rx:csr_write
	signal mm_interconnect_0_sgdma_rx_csr_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:sgdma_rx_csr_writedata -> sgdma_rx:csr_writedata
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                  : std_logic_vector(31 downto 0); -- cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest               : std_logic;                     -- cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess               : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                   : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                      : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                     : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	signal mm_interconnect_0_pb_cpu_to_io_s0_readdata                      : std_logic_vector(31 downto 0); -- pb_cpu_to_io:s0_readdata -> mm_interconnect_0:pb_cpu_to_io_s0_readdata
	signal mm_interconnect_0_pb_cpu_to_io_s0_waitrequest                   : std_logic;                     -- pb_cpu_to_io:s0_waitrequest -> mm_interconnect_0:pb_cpu_to_io_s0_waitrequest
	signal mm_interconnect_0_pb_cpu_to_io_s0_debugaccess                   : std_logic;                     -- mm_interconnect_0:pb_cpu_to_io_s0_debugaccess -> pb_cpu_to_io:s0_debugaccess
	signal mm_interconnect_0_pb_cpu_to_io_s0_address                       : std_logic_vector(9 downto 0);  -- mm_interconnect_0:pb_cpu_to_io_s0_address -> pb_cpu_to_io:s0_address
	signal mm_interconnect_0_pb_cpu_to_io_s0_read                          : std_logic;                     -- mm_interconnect_0:pb_cpu_to_io_s0_read -> pb_cpu_to_io:s0_read
	signal mm_interconnect_0_pb_cpu_to_io_s0_byteenable                    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:pb_cpu_to_io_s0_byteenable -> pb_cpu_to_io:s0_byteenable
	signal mm_interconnect_0_pb_cpu_to_io_s0_readdatavalid                 : std_logic;                     -- pb_cpu_to_io:s0_readdatavalid -> mm_interconnect_0:pb_cpu_to_io_s0_readdatavalid
	signal mm_interconnect_0_pb_cpu_to_io_s0_write                         : std_logic;                     -- mm_interconnect_0:pb_cpu_to_io_s0_write -> pb_cpu_to_io:s0_write
	signal mm_interconnect_0_pb_cpu_to_io_s0_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:pb_cpu_to_io_s0_writedata -> pb_cpu_to_io:s0_writedata
	signal mm_interconnect_0_pb_cpu_to_io_s0_burstcount                    : std_logic_vector(0 downto 0);  -- mm_interconnect_0:pb_cpu_to_io_s0_burstcount -> pb_cpu_to_io:s0_burstcount
	signal mm_interconnect_0_descriptor_memory_s1_chipselect               : std_logic;                     -- mm_interconnect_0:descriptor_memory_s1_chipselect -> descriptor_memory:chipselect
	signal mm_interconnect_0_descriptor_memory_s1_readdata                 : std_logic_vector(31 downto 0); -- descriptor_memory:readdata -> mm_interconnect_0:descriptor_memory_s1_readdata
	signal mm_interconnect_0_descriptor_memory_s1_address                  : std_logic_vector(10 downto 0); -- mm_interconnect_0:descriptor_memory_s1_address -> descriptor_memory:address
	signal mm_interconnect_0_descriptor_memory_s1_byteenable               : std_logic_vector(3 downto 0);  -- mm_interconnect_0:descriptor_memory_s1_byteenable -> descriptor_memory:byteenable
	signal mm_interconnect_0_descriptor_memory_s1_write                    : std_logic;                     -- mm_interconnect_0:descriptor_memory_s1_write -> descriptor_memory:write
	signal mm_interconnect_0_descriptor_memory_s1_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:descriptor_memory_s1_writedata -> descriptor_memory:writedata
	signal mm_interconnect_0_descriptor_memory_s1_clken                    : std_logic;                     -- mm_interconnect_0:descriptor_memory_s1_clken -> descriptor_memory:clken
	signal mm_interconnect_0_onchip_ram_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_chipselect -> onchip_ram:chipselect
	signal mm_interconnect_0_onchip_ram_s1_readdata                        : std_logic_vector(31 downto 0); -- onchip_ram:readdata -> mm_interconnect_0:onchip_ram_s1_readdata
	signal mm_interconnect_0_onchip_ram_s1_address                         : std_logic_vector(18 downto 0); -- mm_interconnect_0:onchip_ram_s1_address -> onchip_ram:address
	signal mm_interconnect_0_onchip_ram_s1_byteenable                      : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_ram_s1_byteenable -> onchip_ram:byteenable
	signal mm_interconnect_0_onchip_ram_s1_write                           : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_write -> onchip_ram:write
	signal mm_interconnect_0_onchip_ram_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_ram_s1_writedata -> onchip_ram:writedata
	signal mm_interconnect_0_onchip_ram_s1_clken                           : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_clken -> onchip_ram:clken
	signal mm_interconnect_0_onchip_ram_s2_chipselect                      : std_logic;                     -- mm_interconnect_0:onchip_ram_s2_chipselect -> onchip_ram:chipselect2
	signal mm_interconnect_0_onchip_ram_s2_readdata                        : std_logic_vector(31 downto 0); -- onchip_ram:readdata2 -> mm_interconnect_0:onchip_ram_s2_readdata
	signal mm_interconnect_0_onchip_ram_s2_address                         : std_logic_vector(18 downto 0); -- mm_interconnect_0:onchip_ram_s2_address -> onchip_ram:address2
	signal mm_interconnect_0_onchip_ram_s2_byteenable                      : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_ram_s2_byteenable -> onchip_ram:byteenable2
	signal mm_interconnect_0_onchip_ram_s2_write                           : std_logic;                     -- mm_interconnect_0:onchip_ram_s2_write -> onchip_ram:write2
	signal mm_interconnect_0_onchip_ram_s2_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_ram_s2_writedata -> onchip_ram:writedata2
	signal mm_interconnect_0_onchip_ram_s2_clken                           : std_logic;                     -- mm_interconnect_0:onchip_ram_s2_clken -> onchip_ram:clken2
	signal pb_cpu_to_io_m0_waitrequest                                     : std_logic;                     -- mm_interconnect_1:pb_cpu_to_io_m0_waitrequest -> pb_cpu_to_io:m0_waitrequest
	signal pb_cpu_to_io_m0_readdata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_1:pb_cpu_to_io_m0_readdata -> pb_cpu_to_io:m0_readdata
	signal pb_cpu_to_io_m0_debugaccess                                     : std_logic;                     -- pb_cpu_to_io:m0_debugaccess -> mm_interconnect_1:pb_cpu_to_io_m0_debugaccess
	signal pb_cpu_to_io_m0_address                                         : std_logic_vector(9 downto 0);  -- pb_cpu_to_io:m0_address -> mm_interconnect_1:pb_cpu_to_io_m0_address
	signal pb_cpu_to_io_m0_read                                            : std_logic;                     -- pb_cpu_to_io:m0_read -> mm_interconnect_1:pb_cpu_to_io_m0_read
	signal pb_cpu_to_io_m0_byteenable                                      : std_logic_vector(3 downto 0);  -- pb_cpu_to_io:m0_byteenable -> mm_interconnect_1:pb_cpu_to_io_m0_byteenable
	signal pb_cpu_to_io_m0_readdatavalid                                   : std_logic;                     -- mm_interconnect_1:pb_cpu_to_io_m0_readdatavalid -> pb_cpu_to_io:m0_readdatavalid
	signal pb_cpu_to_io_m0_writedata                                       : std_logic_vector(31 downto 0); -- pb_cpu_to_io:m0_writedata -> mm_interconnect_1:pb_cpu_to_io_m0_writedata
	signal pb_cpu_to_io_m0_write                                           : std_logic;                     -- pb_cpu_to_io:m0_write -> mm_interconnect_1:pb_cpu_to_io_m0_write
	signal pb_cpu_to_io_m0_burstcount                                      : std_logic_vector(0 downto 0);  -- pb_cpu_to_io:m0_burstcount -> mm_interconnect_1:pb_cpu_to_io_m0_burstcount
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_1_sysid_control_slave_readdata                  : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	signal mm_interconnect_1_sysid_control_slave_address                   : std_logic_vector(0 downto 0);  -- mm_interconnect_1:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_1_sys_clk_timer_s1_chipselect                   : std_logic;                     -- mm_interconnect_1:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	signal mm_interconnect_1_sys_clk_timer_s1_readdata                     : std_logic_vector(15 downto 0); -- sys_clk_timer:readdata -> mm_interconnect_1:sys_clk_timer_s1_readdata
	signal mm_interconnect_1_sys_clk_timer_s1_address                      : std_logic_vector(2 downto 0);  -- mm_interconnect_1:sys_clk_timer_s1_address -> sys_clk_timer:address
	signal mm_interconnect_1_sys_clk_timer_s1_write                        : std_logic;                     -- mm_interconnect_1:sys_clk_timer_s1_write -> mm_interconnect_1_sys_clk_timer_s1_write:in
	signal mm_interconnect_1_sys_clk_timer_s1_writedata                    : std_logic_vector(15 downto 0); -- mm_interconnect_1:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	signal mm_interconnect_1_high_res_timer_s1_chipselect                  : std_logic;                     -- mm_interconnect_1:high_res_timer_s1_chipselect -> high_res_timer:chipselect
	signal mm_interconnect_1_high_res_timer_s1_readdata                    : std_logic_vector(15 downto 0); -- high_res_timer:readdata -> mm_interconnect_1:high_res_timer_s1_readdata
	signal mm_interconnect_1_high_res_timer_s1_address                     : std_logic_vector(2 downto 0);  -- mm_interconnect_1:high_res_timer_s1_address -> high_res_timer:address
	signal mm_interconnect_1_high_res_timer_s1_write                       : std_logic;                     -- mm_interconnect_1:high_res_timer_s1_write -> mm_interconnect_1_high_res_timer_s1_write:in
	signal mm_interconnect_1_high_res_timer_s1_writedata                   : std_logic_vector(15 downto 0); -- mm_interconnect_1:high_res_timer_s1_writedata -> high_res_timer:writedata
	signal irq_mapper_receiver0_irq                                        : std_logic;                     -- sgdma_rx:csr_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                        : std_logic;                     -- sgdma_tx:csr_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                        : std_logic;                     -- sys_clk_timer:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                        : std_logic;                     -- high_res_timer:irq -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                        : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver4_irq
	signal cpu_irq_irq                                                     : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:irq
	signal tse_mac_receive_valid                                           : std_logic;                     -- tse_mac:ff_rx_dval -> avalon_st_adapter:in_0_valid
	signal tse_mac_receive_data                                            : std_logic_vector(31 downto 0); -- tse_mac:ff_rx_data -> avalon_st_adapter:in_0_data
	signal tse_mac_receive_ready                                           : std_logic;                     -- avalon_st_adapter:in_0_ready -> tse_mac:ff_rx_rdy
	signal tse_mac_receive_startofpacket                                   : std_logic;                     -- tse_mac:ff_rx_sop -> avalon_st_adapter:in_0_startofpacket
	signal tse_mac_receive_endofpacket                                     : std_logic;                     -- tse_mac:ff_rx_eop -> avalon_st_adapter:in_0_endofpacket
	signal tse_mac_receive_error                                           : std_logic_vector(5 downto 0);  -- tse_mac:rx_err -> avalon_st_adapter:in_0_error
	signal tse_mac_receive_empty                                           : std_logic_vector(1 downto 0);  -- tse_mac:ff_rx_mod -> avalon_st_adapter:in_0_empty
	signal avalon_st_adapter_out_0_valid                                   : std_logic;                     -- avalon_st_adapter:out_0_valid -> sgdma_rx:in_valid
	signal avalon_st_adapter_out_0_data                                    : std_logic_vector(31 downto 0); -- avalon_st_adapter:out_0_data -> sgdma_rx:in_data
	signal avalon_st_adapter_out_0_ready                                   : std_logic;                     -- sgdma_rx:in_ready -> avalon_st_adapter:out_0_ready
	signal avalon_st_adapter_out_0_startofpacket                           : std_logic;                     -- avalon_st_adapter:out_0_startofpacket -> sgdma_rx:in_startofpacket
	signal avalon_st_adapter_out_0_endofpacket                             : std_logic;                     -- avalon_st_adapter:out_0_endofpacket -> sgdma_rx:in_endofpacket
	signal avalon_st_adapter_out_0_error                                   : std_logic_vector(5 downto 0);  -- avalon_st_adapter:out_0_error -> sgdma_rx:in_error
	signal avalon_st_adapter_out_0_empty                                   : std_logic_vector(1 downto 0);  -- avalon_st_adapter:out_0_empty -> sgdma_rx:in_empty
	signal rst_controller_reset_out_reset                                  : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, mm_interconnect_1:pb_cpu_to_io_reset_reset_bridge_in_reset_reset, pb_cpu_to_io:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                              : std_logic;                     -- rst_controller:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	signal cpu_debug_reset_request_reset                                   : std_logic;                     -- cpu:debug_reset_request -> rst_controller:reset_in1
	signal rst_controller_001_reset_out_reset                              : std_logic;                     -- rst_controller_001:reset_out -> [avalon_st_adapter:in_rst_0_reset, descriptor_memory:reset, mm_interconnect_0:sgdma_rx_reset_reset_bridge_in_reset_reset, mm_interconnect_1:jtag_uart_0_reset_reset_bridge_in_reset_reset, onchip_ram:reset, onchip_ram:reset2, rst_controller_001_reset_out_reset:in, rst_translator_001:in_reset, tse_mac:reset]
	signal rst_controller_001_reset_out_reset_req                          : std_logic;                     -- rst_controller_001:reset_req -> [descriptor_memory:reset_req, onchip_ram:reset_req, onchip_ram:reset_req2, rst_translator_001:reset_req_in]
	signal rst_controller_002_reset_out_reset                              : std_logic;                     -- rst_controller_002:reset_out -> [mm_interconnect_0:mem_if_lpddr2_emif_0_avl_0_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:mem_if_lpddr2_emif_0_mp_cmd_reset_n_0_reset_bridge_in_reset_reset]
	signal merged_resets_in_reset_reset_n_ports_inv                        : std_logic;                     -- merged_resets_in_reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller:reset_in2, rst_controller_001:reset_in0, rst_controller_001:reset_in1, rst_controller_002:reset_in0]
	signal mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_inv                : std_logic;                     -- mem_if_lpddr2_emif_0_avl_0_waitrequest:inv -> mm_interconnect_0:mem_if_lpddr2_emif_0_avl_0_waitrequest
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_1_sys_clk_timer_s1_write_ports_inv              : std_logic;                     -- mm_interconnect_1_sys_clk_timer_s1_write:inv -> sys_clk_timer:write_n
	signal mm_interconnect_1_high_res_timer_s1_write_ports_inv             : std_logic;                     -- mm_interconnect_1_high_res_timer_s1_write:inv -> high_res_timer:write_n
	signal rst_controller_reset_out_reset_ports_inv                        : std_logic;                     -- rst_controller_reset_out_reset:inv -> cpu:reset_n
	signal rst_controller_001_reset_out_reset_ports_inv                    : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [high_res_timer:reset_n, jtag_uart_0:rst_n, sgdma_rx:system_reset_n, sgdma_tx:system_reset_n, sys_clk_timer:reset_n, sysid:reset_n]

begin

	cpu : component Nios_CPU_qsys_cpu
		port map (
			clk                                 => clk_clk,                                           --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,          --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => cpu_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	descriptor_memory : component Nios_CPU_qsys_descriptor_memory
		port map (
			clk        => clk_clk,                                           --   clk1.clk
			address    => mm_interconnect_0_descriptor_memory_s1_address,    --     s1.address
			clken      => mm_interconnect_0_descriptor_memory_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_descriptor_memory_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_descriptor_memory_s1_write,      --       .write
			readdata   => mm_interconnect_0_descriptor_memory_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_descriptor_memory_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_descriptor_memory_s1_byteenable, --       .byteenable
			reset      => rst_controller_001_reset_out_reset,                -- reset1.reset
			reset_req  => rst_controller_001_reset_out_reset_req,            --       .reset_req
			freeze     => '0'                                                -- (terminated)
		);

	high_res_timer : component Nios_CPU_qsys_high_res_timer
		port map (
			clk        => clk_clk,                                             --   clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,        -- reset.reset_n
			address    => mm_interconnect_1_high_res_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_1_high_res_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_1_high_res_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_1_high_res_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_1_high_res_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver3_irq                             --   irq.irq
		);

	jtag_uart_0 : component Nios_CPU_qsys_jtag_uart_0
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                    --             reset.reset_n
			av_chipselect  => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver4_irq                                         --               irq.irq
		);

	mem_if_lpddr2_emif_0 : component Nios_CPU_qsys_mem_if_lpddr2_emif_0
		port map (
			pll_ref_clk                => clk_clk,                                                         --        pll_ref_clk.clk
			global_reset_n             => merged_resets_in_reset_reset_n,                                  --       global_reset.reset_n
			soft_reset_n               => merged_resets_in_reset_reset_n,                                  --         soft_reset.reset_n
			afi_clk                    => mem_if_lpddr2_emif_0_afi_clk_clk,                                --            afi_clk.clk
			afi_half_clk               => open,                                                            --       afi_half_clk.clk
			afi_reset_n                => open,                                                            --          afi_reset.reset_n
			afi_reset_export_n         => open,                                                            --   afi_reset_export.reset_n
			mem_ca                     => memory_mem_ca,                                                   --             memory.mem_ca
			mem_ck                     => memory_mem_ck,                                                   --                   .mem_ck
			mem_ck_n                   => memory_mem_ck_n,                                                 --                   .mem_ck_n
			mem_cke                    => memory_mem_cke,                                                  --                   .mem_cke
			mem_cs_n                   => memory_mem_cs_n,                                                 --                   .mem_cs_n
			mem_dm                     => memory_mem_dm,                                                   --                   .mem_dm
			mem_dq                     => memory_mem_dq,                                                   --                   .mem_dq
			mem_dqs                    => memory_mem_dqs,                                                  --                   .mem_dqs
			mem_dqs_n                  => memory_mem_dqs_n,                                                --                   .mem_dqs_n
			avl_ready_0                => mem_if_lpddr2_emif_0_avl_0_waitrequest,                          --              avl_0.waitrequest_n
			avl_burstbegin_0           => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_beginbursttransfer, --                   .beginbursttransfer
			avl_addr_0                 => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_address,            --                   .address
			avl_rdata_valid_0          => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_readdatavalid,      --                   .readdatavalid
			avl_rdata_0                => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_readdata,           --                   .readdata
			avl_wdata_0                => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_writedata,          --                   .writedata
			avl_be_0                   => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_byteenable,         --                   .byteenable
			avl_read_req_0             => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_read,               --                   .read
			avl_write_req_0            => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_write,              --                   .write
			avl_size_0                 => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_burstcount,         --                   .burstcount
			mp_cmd_clk_0_clk           => mem_if_lpddr2_emif_0_afi_clk_clk,                                --       mp_cmd_clk_0.clk
			mp_cmd_reset_n_0_reset_n   => merged_resets_in_reset_reset_n,                                  --   mp_cmd_reset_n_0.reset_n
			mp_rfifo_clk_0_clk         => mem_if_lpddr2_emif_0_afi_clk_clk,                                --     mp_rfifo_clk_0.clk
			mp_rfifo_reset_n_0_reset_n => merged_resets_in_reset_reset_n,                                  -- mp_rfifo_reset_n_0.reset_n
			mp_wfifo_clk_0_clk         => mem_if_lpddr2_emif_0_afi_clk_clk,                                --     mp_wfifo_clk_0.clk
			mp_wfifo_reset_n_0_reset_n => merged_resets_in_reset_reset_n,                                  -- mp_wfifo_reset_n_0.reset_n
			local_init_done            => mem_if_lpddr2_emif_0_status_local_init_done,                     --             status.local_init_done
			local_cal_success          => mem_if_lpddr2_emif_0_status_local_cal_success,                   --                   .local_cal_success
			local_cal_fail             => mem_if_lpddr2_emif_0_status_local_cal_fail,                      --                   .local_cal_fail
			oct_rzqin                  => oct_rzqin,                                                       --                oct.rzqin
			pll_mem_clk                => mem_if_lpddr2_emif_0_pll_sharing_pll_mem_clk,                    --        pll_sharing.pll_mem_clk
			pll_write_clk              => mem_if_lpddr2_emif_0_pll_sharing_pll_write_clk,                  --                   .pll_write_clk
			pll_locked                 => mem_if_lpddr2_emif_0_pll_sharing_pll_locked,                     --                   .pll_locked
			pll_write_clk_pre_phy_clk  => mem_if_lpddr2_emif_0_pll_sharing_pll_write_clk_pre_phy_clk,      --                   .pll_write_clk_pre_phy_clk
			pll_addr_cmd_clk           => mem_if_lpddr2_emif_0_pll_sharing_pll_addr_cmd_clk,               --                   .pll_addr_cmd_clk
			pll_avl_clk                => mem_if_lpddr2_emif_0_pll_sharing_pll_avl_clk,                    --                   .pll_avl_clk
			pll_config_clk             => mem_if_lpddr2_emif_0_pll_sharing_pll_config_clk,                 --                   .pll_config_clk
			pll_mem_phy_clk            => mem_if_lpddr2_emif_0_pll_sharing_pll_mem_phy_clk,                --                   .pll_mem_phy_clk
			afi_phy_clk                => mem_if_lpddr2_emif_0_pll_sharing_afi_phy_clk,                    --                   .afi_phy_clk
			pll_avl_phy_clk            => mem_if_lpddr2_emif_0_pll_sharing_pll_avl_phy_clk                 --                   .pll_avl_phy_clk
		);

	onchip_ram : component Nios_CPU_qsys_onchip_ram
		port map (
			clk         => clk_clk,                                    --   clk1.clk
			address     => mm_interconnect_0_onchip_ram_s1_address,    --     s1.address
			clken       => mm_interconnect_0_onchip_ram_s1_clken,      --       .clken
			chipselect  => mm_interconnect_0_onchip_ram_s1_chipselect, --       .chipselect
			write       => mm_interconnect_0_onchip_ram_s1_write,      --       .write
			readdata    => mm_interconnect_0_onchip_ram_s1_readdata,   --       .readdata
			writedata   => mm_interconnect_0_onchip_ram_s1_writedata,  --       .writedata
			byteenable  => mm_interconnect_0_onchip_ram_s1_byteenable, --       .byteenable
			reset       => rst_controller_001_reset_out_reset,         -- reset1.reset
			reset_req   => rst_controller_001_reset_out_reset_req,     --       .reset_req
			address2    => mm_interconnect_0_onchip_ram_s2_address,    --     s2.address
			chipselect2 => mm_interconnect_0_onchip_ram_s2_chipselect, --       .chipselect
			clken2      => mm_interconnect_0_onchip_ram_s2_clken,      --       .clken
			write2      => mm_interconnect_0_onchip_ram_s2_write,      --       .write
			readdata2   => mm_interconnect_0_onchip_ram_s2_readdata,   --       .readdata
			writedata2  => mm_interconnect_0_onchip_ram_s2_writedata,  --       .writedata
			byteenable2 => mm_interconnect_0_onchip_ram_s2_byteenable, --       .byteenable
			clk2        => clk_clk,                                    --   clk2.clk
			reset2      => rst_controller_001_reset_out_reset,         -- reset2.reset
			reset_req2  => rst_controller_001_reset_out_reset_req,     --       .reset_req
			freeze      => '0'                                         -- (terminated)
		);

	pb_cpu_to_io : component altera_avalon_mm_bridge
		generic map (
			DATA_WIDTH        => 32,
			SYMBOL_WIDTH      => 8,
			HDL_ADDR_WIDTH    => 10,
			BURSTCOUNT_WIDTH  => 1,
			PIPELINE_COMMAND  => 1,
			PIPELINE_RESPONSE => 1
		)
		port map (
			clk              => clk_clk,                                         --   clk.clk
			reset            => rst_controller_reset_out_reset,                  -- reset.reset
			s0_waitrequest   => mm_interconnect_0_pb_cpu_to_io_s0_waitrequest,   --    s0.waitrequest
			s0_readdata      => mm_interconnect_0_pb_cpu_to_io_s0_readdata,      --      .readdata
			s0_readdatavalid => mm_interconnect_0_pb_cpu_to_io_s0_readdatavalid, --      .readdatavalid
			s0_burstcount    => mm_interconnect_0_pb_cpu_to_io_s0_burstcount,    --      .burstcount
			s0_writedata     => mm_interconnect_0_pb_cpu_to_io_s0_writedata,     --      .writedata
			s0_address       => mm_interconnect_0_pb_cpu_to_io_s0_address,       --      .address
			s0_write         => mm_interconnect_0_pb_cpu_to_io_s0_write,         --      .write
			s0_read          => mm_interconnect_0_pb_cpu_to_io_s0_read,          --      .read
			s0_byteenable    => mm_interconnect_0_pb_cpu_to_io_s0_byteenable,    --      .byteenable
			s0_debugaccess   => mm_interconnect_0_pb_cpu_to_io_s0_debugaccess,   --      .debugaccess
			m0_waitrequest   => pb_cpu_to_io_m0_waitrequest,                     --    m0.waitrequest
			m0_readdata      => pb_cpu_to_io_m0_readdata,                        --      .readdata
			m0_readdatavalid => pb_cpu_to_io_m0_readdatavalid,                   --      .readdatavalid
			m0_burstcount    => pb_cpu_to_io_m0_burstcount,                      --      .burstcount
			m0_writedata     => pb_cpu_to_io_m0_writedata,                       --      .writedata
			m0_address       => pb_cpu_to_io_m0_address,                         --      .address
			m0_write         => pb_cpu_to_io_m0_write,                           --      .write
			m0_read          => pb_cpu_to_io_m0_read,                            --      .read
			m0_byteenable    => pb_cpu_to_io_m0_byteenable,                      --      .byteenable
			m0_debugaccess   => pb_cpu_to_io_m0_debugaccess,                     --      .debugaccess
			s0_response      => open,                                            -- (terminated)
			m0_response      => "00"                                             -- (terminated)
		);

	sgdma_rx : component Nios_CPU_qsys_sgdma_rx
		port map (
			clk                           => clk_clk,                                      --              clk.clk
			system_reset_n                => rst_controller_001_reset_out_reset_ports_inv, --            reset.reset_n
			csr_chipselect                => mm_interconnect_0_sgdma_rx_csr_chipselect,    --              csr.chipselect
			csr_address                   => mm_interconnect_0_sgdma_rx_csr_address,       --                 .address
			csr_read                      => mm_interconnect_0_sgdma_rx_csr_read,          --                 .read
			csr_write                     => mm_interconnect_0_sgdma_rx_csr_write,         --                 .write
			csr_writedata                 => mm_interconnect_0_sgdma_rx_csr_writedata,     --                 .writedata
			csr_readdata                  => mm_interconnect_0_sgdma_rx_csr_readdata,      --                 .readdata
			descriptor_read_readdata      => sgdma_rx_descriptor_read_readdata,            --  descriptor_read.readdata
			descriptor_read_readdatavalid => sgdma_rx_descriptor_read_readdatavalid,       --                 .readdatavalid
			descriptor_read_waitrequest   => sgdma_rx_descriptor_read_waitrequest,         --                 .waitrequest
			descriptor_read_address       => sgdma_rx_descriptor_read_address,             --                 .address
			descriptor_read_read          => sgdma_rx_descriptor_read_read,                --                 .read
			descriptor_write_waitrequest  => sgdma_rx_descriptor_write_waitrequest,        -- descriptor_write.waitrequest
			descriptor_write_address      => sgdma_rx_descriptor_write_address,            --                 .address
			descriptor_write_write        => sgdma_rx_descriptor_write_write,              --                 .write
			descriptor_write_writedata    => sgdma_rx_descriptor_write_writedata,          --                 .writedata
			csr_irq                       => irq_mapper_receiver0_irq,                     --          csr_irq.irq
			in_startofpacket              => avalon_st_adapter_out_0_startofpacket,        --               in.startofpacket
			in_endofpacket                => avalon_st_adapter_out_0_endofpacket,          --                 .endofpacket
			in_data                       => avalon_st_adapter_out_0_data,                 --                 .data
			in_valid                      => avalon_st_adapter_out_0_valid,                --                 .valid
			in_ready                      => avalon_st_adapter_out_0_ready,                --                 .ready
			in_empty                      => avalon_st_adapter_out_0_empty,                --                 .empty
			in_error                      => avalon_st_adapter_out_0_error,                --                 .error
			m_write_waitrequest           => sgdma_rx_m_write_waitrequest,                 --          m_write.waitrequest
			m_write_address               => sgdma_rx_m_write_address,                     --                 .address
			m_write_write                 => sgdma_rx_m_write_write,                       --                 .write
			m_write_writedata             => sgdma_rx_m_write_writedata,                   --                 .writedata
			m_write_byteenable            => sgdma_rx_m_write_byteenable                   --                 .byteenable
		);

	sgdma_tx : component Nios_CPU_qsys_sgdma_tx
		port map (
			clk                           => clk_clk,                                      --              clk.clk
			system_reset_n                => rst_controller_001_reset_out_reset_ports_inv, --            reset.reset_n
			csr_chipselect                => mm_interconnect_0_sgdma_tx_csr_chipselect,    --              csr.chipselect
			csr_address                   => mm_interconnect_0_sgdma_tx_csr_address,       --                 .address
			csr_read                      => mm_interconnect_0_sgdma_tx_csr_read,          --                 .read
			csr_write                     => mm_interconnect_0_sgdma_tx_csr_write,         --                 .write
			csr_writedata                 => mm_interconnect_0_sgdma_tx_csr_writedata,     --                 .writedata
			csr_readdata                  => mm_interconnect_0_sgdma_tx_csr_readdata,      --                 .readdata
			descriptor_read_readdata      => sgdma_tx_descriptor_read_readdata,            --  descriptor_read.readdata
			descriptor_read_readdatavalid => sgdma_tx_descriptor_read_readdatavalid,       --                 .readdatavalid
			descriptor_read_waitrequest   => sgdma_tx_descriptor_read_waitrequest,         --                 .waitrequest
			descriptor_read_address       => sgdma_tx_descriptor_read_address,             --                 .address
			descriptor_read_read          => sgdma_tx_descriptor_read_read,                --                 .read
			descriptor_write_waitrequest  => sgdma_tx_descriptor_write_waitrequest,        -- descriptor_write.waitrequest
			descriptor_write_address      => sgdma_tx_descriptor_write_address,            --                 .address
			descriptor_write_write        => sgdma_tx_descriptor_write_write,              --                 .write
			descriptor_write_writedata    => sgdma_tx_descriptor_write_writedata,          --                 .writedata
			csr_irq                       => irq_mapper_receiver1_irq,                     --          csr_irq.irq
			m_read_readdata               => sgdma_tx_m_read_readdata,                     --           m_read.readdata
			m_read_readdatavalid          => sgdma_tx_m_read_readdatavalid,                --                 .readdatavalid
			m_read_waitrequest            => sgdma_tx_m_read_waitrequest,                  --                 .waitrequest
			m_read_address                => sgdma_tx_m_read_address,                      --                 .address
			m_read_read                   => sgdma_tx_m_read_read,                         --                 .read
			out_data                      => sgdma_tx_out_data,                            --              out.data
			out_valid                     => sgdma_tx_out_valid,                           --                 .valid
			out_ready                     => sgdma_tx_out_ready,                           --                 .ready
			out_endofpacket               => sgdma_tx_out_endofpacket,                     --                 .endofpacket
			out_startofpacket             => sgdma_tx_out_startofpacket,                   --                 .startofpacket
			out_empty                     => sgdma_tx_out_empty,                           --                 .empty
			out_error                     => sgdma_tx_out_error                            --                 .error
		);

	sys_clk_timer : component Nios_CPU_qsys_sys_clk_timer
		port map (
			clk        => clk_clk,                                            --   clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,       -- reset.reset_n
			address    => mm_interconnect_1_sys_clk_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_1_sys_clk_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_1_sys_clk_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_1_sys_clk_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_1_sys_clk_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver2_irq                            --   irq.irq
		);

	sysid : component Nios_CPU_qsys_sysid
		port map (
			clock    => clk_clk,                                          --           clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,     --         reset.reset_n
			readdata => mm_interconnect_1_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_1_sysid_control_slave_address(0)  --              .address
		);

	tse_mac : component Nios_CPU_qsys_tse_mac
		port map (
			clk           => clk_clk,                                            -- control_port_clock_connection.clk
			reset         => rst_controller_001_reset_out_reset,                 --              reset_connection.reset
			reg_addr      => mm_interconnect_0_tse_mac_control_port_address,     --                  control_port.address
			reg_data_out  => mm_interconnect_0_tse_mac_control_port_readdata,    --                              .readdata
			reg_rd        => mm_interconnect_0_tse_mac_control_port_read,        --                              .read
			reg_data_in   => mm_interconnect_0_tse_mac_control_port_writedata,   --                              .writedata
			reg_wr        => mm_interconnect_0_tse_mac_control_port_write,       --                              .write
			reg_busy      => mm_interconnect_0_tse_mac_control_port_waitrequest, --                              .waitrequest
			tx_clk        => tse_mac_pcs_mac_tx_clock_connection_clk,            --   pcs_mac_tx_clock_connection.clk
			rx_clk        => tse_mac_pcs_mac_rx_clock_connection_clk,            --   pcs_mac_rx_clock_connection.clk
			set_10        => tse_mac_mac_status_connection_set_10,               --         mac_status_connection.set_10
			set_1000      => tse_mac_mac_status_connection_set_1000,             --                              .set_1000
			eth_mode      => tse_mac_mac_status_connection_eth_mode,             --                              .eth_mode
			ena_10        => tse_mac_mac_status_connection_ena_10,               --                              .ena_10
			gm_rx_d       => tse_mac_mac_gmii_connection_gmii_rx_d,              --           mac_gmii_connection.gmii_rx_d
			gm_rx_dv      => tse_mac_mac_gmii_connection_gmii_rx_dv,             --                              .gmii_rx_dv
			gm_rx_err     => tse_mac_mac_gmii_connection_gmii_rx_err,            --                              .gmii_rx_err
			gm_tx_d       => tse_mac_mac_gmii_connection_gmii_tx_d,              --                              .gmii_tx_d
			gm_tx_en      => tse_mac_mac_gmii_connection_gmii_tx_en,             --                              .gmii_tx_en
			gm_tx_err     => tse_mac_mac_gmii_connection_gmii_tx_err,            --                              .gmii_tx_err
			m_rx_d        => tse_mac_mac_mii_connection_mii_rx_d,                --            mac_mii_connection.mii_rx_d
			m_rx_en       => tse_mac_mac_mii_connection_mii_rx_dv,               --                              .mii_rx_dv
			m_rx_err      => tse_mac_mac_mii_connection_mii_rx_err,              --                              .mii_rx_err
			m_tx_d        => tse_mac_mac_mii_connection_mii_tx_d,                --                              .mii_tx_d
			m_tx_en       => tse_mac_mac_mii_connection_mii_tx_en,               --                              .mii_tx_en
			m_tx_err      => tse_mac_mac_mii_connection_mii_tx_err,              --                              .mii_tx_err
			m_rx_crs      => tse_mac_mac_mii_connection_mii_crs,                 --                              .mii_crs
			m_rx_col      => tse_mac_mac_mii_connection_mii_col,                 --                              .mii_col
			ff_rx_clk     => clk_clk,                                            --      receive_clock_connection.clk
			ff_tx_clk     => clk_clk,                                            --     transmit_clock_connection.clk
			ff_rx_data    => tse_mac_receive_data,                               --                       receive.data
			ff_rx_eop     => tse_mac_receive_endofpacket,                        --                              .endofpacket
			rx_err        => tse_mac_receive_error,                              --                              .error
			ff_rx_mod     => tse_mac_receive_empty,                              --                              .empty
			ff_rx_rdy     => tse_mac_receive_ready,                              --                              .ready
			ff_rx_sop     => tse_mac_receive_startofpacket,                      --                              .startofpacket
			ff_rx_dval    => tse_mac_receive_valid,                              --                              .valid
			ff_tx_data    => sgdma_tx_out_data,                                  --                      transmit.data
			ff_tx_eop     => sgdma_tx_out_endofpacket,                           --                              .endofpacket
			ff_tx_err     => sgdma_tx_out_error,                                 --                              .error
			ff_tx_mod     => sgdma_tx_out_empty,                                 --                              .empty
			ff_tx_rdy     => sgdma_tx_out_ready,                                 --                              .ready
			ff_tx_sop     => sgdma_tx_out_startofpacket,                         --                              .startofpacket
			ff_tx_wren    => sgdma_tx_out_valid,                                 --                              .valid
			mdc           => tse_mac_mac_mdio_connection_mdc,                    --           mac_mdio_connection.mdc
			mdio_in       => tse_mac_mac_mdio_connection_mdio_in,                --                              .mdio_in
			mdio_out      => tse_mac_mac_mdio_connection_mdio_out,               --                              .mdio_out
			mdio_oen      => tse_mac_mac_mdio_connection_mdio_oen,               --                              .mdio_oen
			xon_gen       => tse_mac_mac_misc_connection_xon_gen,                --           mac_misc_connection.xon_gen
			xoff_gen      => tse_mac_mac_misc_connection_xoff_gen,               --                              .xoff_gen
			ff_tx_crc_fwd => tse_mac_mac_misc_connection_ff_tx_crc_fwd,          --                              .ff_tx_crc_fwd
			ff_tx_septy   => tse_mac_mac_misc_connection_ff_tx_septy,            --                              .ff_tx_septy
			tx_ff_uflow   => tse_mac_mac_misc_connection_tx_ff_uflow,            --                              .tx_ff_uflow
			ff_tx_a_full  => tse_mac_mac_misc_connection_ff_tx_a_full,           --                              .ff_tx_a_full
			ff_tx_a_empty => tse_mac_mac_misc_connection_ff_tx_a_empty,          --                              .ff_tx_a_empty
			rx_err_stat   => tse_mac_mac_misc_connection_rx_err_stat,            --                              .rx_err_stat
			rx_frm_type   => tse_mac_mac_misc_connection_rx_frm_type,            --                              .rx_frm_type
			ff_rx_dsav    => tse_mac_mac_misc_connection_ff_rx_dsav,             --                              .ff_rx_dsav
			ff_rx_a_full  => tse_mac_mac_misc_connection_ff_rx_a_full,           --                              .ff_rx_a_full
			ff_rx_a_empty => tse_mac_mac_misc_connection_ff_rx_a_empty           --                              .ff_rx_a_empty
		);

	mm_interconnect_0 : component Nios_CPU_qsys_mm_interconnect_0
		port map (
			clkin_50_clk_clk                                                        => clk_clk,                                                         --                                                      clkin_50_clk.clk
			mem_if_lpddr2_emif_0_afi_clk_clk                                        => mem_if_lpddr2_emif_0_afi_clk_clk,                                --                                      mem_if_lpddr2_emif_0_afi_clk.clk
			cpu_reset_reset_bridge_in_reset_reset                                   => rst_controller_reset_out_reset,                                  --                                   cpu_reset_reset_bridge_in_reset.reset
			mem_if_lpddr2_emif_0_avl_0_translator_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                              -- mem_if_lpddr2_emif_0_avl_0_translator_reset_reset_bridge_in_reset.reset
			mem_if_lpddr2_emif_0_mp_cmd_reset_n_0_reset_bridge_in_reset_reset       => rst_controller_002_reset_out_reset,                              --       mem_if_lpddr2_emif_0_mp_cmd_reset_n_0_reset_bridge_in_reset.reset
			sgdma_rx_reset_reset_bridge_in_reset_reset                              => rst_controller_001_reset_out_reset,                              --                              sgdma_rx_reset_reset_bridge_in_reset.reset
			cpu_data_master_address                                                 => cpu_data_master_address,                                         --                                                   cpu_data_master.address
			cpu_data_master_waitrequest                                             => cpu_data_master_waitrequest,                                     --                                                                  .waitrequest
			cpu_data_master_byteenable                                              => cpu_data_master_byteenable,                                      --                                                                  .byteenable
			cpu_data_master_read                                                    => cpu_data_master_read,                                            --                                                                  .read
			cpu_data_master_readdata                                                => cpu_data_master_readdata,                                        --                                                                  .readdata
			cpu_data_master_readdatavalid                                           => cpu_data_master_readdatavalid,                                   --                                                                  .readdatavalid
			cpu_data_master_write                                                   => cpu_data_master_write,                                           --                                                                  .write
			cpu_data_master_writedata                                               => cpu_data_master_writedata,                                       --                                                                  .writedata
			cpu_data_master_debugaccess                                             => cpu_data_master_debugaccess,                                     --                                                                  .debugaccess
			cpu_instruction_master_address                                          => cpu_instruction_master_address,                                  --                                            cpu_instruction_master.address
			cpu_instruction_master_waitrequest                                      => cpu_instruction_master_waitrequest,                              --                                                                  .waitrequest
			cpu_instruction_master_read                                             => cpu_instruction_master_read,                                     --                                                                  .read
			cpu_instruction_master_readdata                                         => cpu_instruction_master_readdata,                                 --                                                                  .readdata
			cpu_instruction_master_readdatavalid                                    => cpu_instruction_master_readdatavalid,                            --                                                                  .readdatavalid
			sgdma_rx_descriptor_read_address                                        => sgdma_rx_descriptor_read_address,                                --                                          sgdma_rx_descriptor_read.address
			sgdma_rx_descriptor_read_waitrequest                                    => sgdma_rx_descriptor_read_waitrequest,                            --                                                                  .waitrequest
			sgdma_rx_descriptor_read_read                                           => sgdma_rx_descriptor_read_read,                                   --                                                                  .read
			sgdma_rx_descriptor_read_readdata                                       => sgdma_rx_descriptor_read_readdata,                               --                                                                  .readdata
			sgdma_rx_descriptor_read_readdatavalid                                  => sgdma_rx_descriptor_read_readdatavalid,                          --                                                                  .readdatavalid
			sgdma_rx_descriptor_write_address                                       => sgdma_rx_descriptor_write_address,                               --                                         sgdma_rx_descriptor_write.address
			sgdma_rx_descriptor_write_waitrequest                                   => sgdma_rx_descriptor_write_waitrequest,                           --                                                                  .waitrequest
			sgdma_rx_descriptor_write_write                                         => sgdma_rx_descriptor_write_write,                                 --                                                                  .write
			sgdma_rx_descriptor_write_writedata                                     => sgdma_rx_descriptor_write_writedata,                             --                                                                  .writedata
			sgdma_rx_m_write_address                                                => sgdma_rx_m_write_address,                                        --                                                  sgdma_rx_m_write.address
			sgdma_rx_m_write_waitrequest                                            => sgdma_rx_m_write_waitrequest,                                    --                                                                  .waitrequest
			sgdma_rx_m_write_byteenable                                             => sgdma_rx_m_write_byteenable,                                     --                                                                  .byteenable
			sgdma_rx_m_write_write                                                  => sgdma_rx_m_write_write,                                          --                                                                  .write
			sgdma_rx_m_write_writedata                                              => sgdma_rx_m_write_writedata,                                      --                                                                  .writedata
			sgdma_tx_descriptor_read_address                                        => sgdma_tx_descriptor_read_address,                                --                                          sgdma_tx_descriptor_read.address
			sgdma_tx_descriptor_read_waitrequest                                    => sgdma_tx_descriptor_read_waitrequest,                            --                                                                  .waitrequest
			sgdma_tx_descriptor_read_read                                           => sgdma_tx_descriptor_read_read,                                   --                                                                  .read
			sgdma_tx_descriptor_read_readdata                                       => sgdma_tx_descriptor_read_readdata,                               --                                                                  .readdata
			sgdma_tx_descriptor_read_readdatavalid                                  => sgdma_tx_descriptor_read_readdatavalid,                          --                                                                  .readdatavalid
			sgdma_tx_descriptor_write_address                                       => sgdma_tx_descriptor_write_address,                               --                                         sgdma_tx_descriptor_write.address
			sgdma_tx_descriptor_write_waitrequest                                   => sgdma_tx_descriptor_write_waitrequest,                           --                                                                  .waitrequest
			sgdma_tx_descriptor_write_write                                         => sgdma_tx_descriptor_write_write,                                 --                                                                  .write
			sgdma_tx_descriptor_write_writedata                                     => sgdma_tx_descriptor_write_writedata,                             --                                                                  .writedata
			sgdma_tx_m_read_address                                                 => sgdma_tx_m_read_address,                                         --                                                   sgdma_tx_m_read.address
			sgdma_tx_m_read_waitrequest                                             => sgdma_tx_m_read_waitrequest,                                     --                                                                  .waitrequest
			sgdma_tx_m_read_read                                                    => sgdma_tx_m_read_read,                                            --                                                                  .read
			sgdma_tx_m_read_readdata                                                => sgdma_tx_m_read_readdata,                                        --                                                                  .readdata
			sgdma_tx_m_read_readdatavalid                                           => sgdma_tx_m_read_readdatavalid,                                   --                                                                  .readdatavalid
			cpu_debug_mem_slave_address                                             => mm_interconnect_0_cpu_debug_mem_slave_address,                   --                                               cpu_debug_mem_slave.address
			cpu_debug_mem_slave_write                                               => mm_interconnect_0_cpu_debug_mem_slave_write,                     --                                                                  .write
			cpu_debug_mem_slave_read                                                => mm_interconnect_0_cpu_debug_mem_slave_read,                      --                                                                  .read
			cpu_debug_mem_slave_readdata                                            => mm_interconnect_0_cpu_debug_mem_slave_readdata,                  --                                                                  .readdata
			cpu_debug_mem_slave_writedata                                           => mm_interconnect_0_cpu_debug_mem_slave_writedata,                 --                                                                  .writedata
			cpu_debug_mem_slave_byteenable                                          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,                --                                                                  .byteenable
			cpu_debug_mem_slave_waitrequest                                         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,               --                                                                  .waitrequest
			cpu_debug_mem_slave_debugaccess                                         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,               --                                                                  .debugaccess
			descriptor_memory_s1_address                                            => mm_interconnect_0_descriptor_memory_s1_address,                  --                                              descriptor_memory_s1.address
			descriptor_memory_s1_write                                              => mm_interconnect_0_descriptor_memory_s1_write,                    --                                                                  .write
			descriptor_memory_s1_readdata                                           => mm_interconnect_0_descriptor_memory_s1_readdata,                 --                                                                  .readdata
			descriptor_memory_s1_writedata                                          => mm_interconnect_0_descriptor_memory_s1_writedata,                --                                                                  .writedata
			descriptor_memory_s1_byteenable                                         => mm_interconnect_0_descriptor_memory_s1_byteenable,               --                                                                  .byteenable
			descriptor_memory_s1_chipselect                                         => mm_interconnect_0_descriptor_memory_s1_chipselect,               --                                                                  .chipselect
			descriptor_memory_s1_clken                                              => mm_interconnect_0_descriptor_memory_s1_clken,                    --                                                                  .clken
			mem_if_lpddr2_emif_0_avl_0_address                                      => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_address,            --                                        mem_if_lpddr2_emif_0_avl_0.address
			mem_if_lpddr2_emif_0_avl_0_write                                        => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_write,              --                                                                  .write
			mem_if_lpddr2_emif_0_avl_0_read                                         => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_read,               --                                                                  .read
			mem_if_lpddr2_emif_0_avl_0_readdata                                     => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_readdata,           --                                                                  .readdata
			mem_if_lpddr2_emif_0_avl_0_writedata                                    => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_writedata,          --                                                                  .writedata
			mem_if_lpddr2_emif_0_avl_0_beginbursttransfer                           => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_beginbursttransfer, --                                                                  .beginbursttransfer
			mem_if_lpddr2_emif_0_avl_0_burstcount                                   => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_burstcount,         --                                                                  .burstcount
			mem_if_lpddr2_emif_0_avl_0_byteenable                                   => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_byteenable,         --                                                                  .byteenable
			mem_if_lpddr2_emif_0_avl_0_readdatavalid                                => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_readdatavalid,      --                                                                  .readdatavalid
			mem_if_lpddr2_emif_0_avl_0_waitrequest                                  => mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_inv,                --                                                                  .waitrequest
			onchip_ram_s1_address                                                   => mm_interconnect_0_onchip_ram_s1_address,                         --                                                     onchip_ram_s1.address
			onchip_ram_s1_write                                                     => mm_interconnect_0_onchip_ram_s1_write,                           --                                                                  .write
			onchip_ram_s1_readdata                                                  => mm_interconnect_0_onchip_ram_s1_readdata,                        --                                                                  .readdata
			onchip_ram_s1_writedata                                                 => mm_interconnect_0_onchip_ram_s1_writedata,                       --                                                                  .writedata
			onchip_ram_s1_byteenable                                                => mm_interconnect_0_onchip_ram_s1_byteenable,                      --                                                                  .byteenable
			onchip_ram_s1_chipselect                                                => mm_interconnect_0_onchip_ram_s1_chipselect,                      --                                                                  .chipselect
			onchip_ram_s1_clken                                                     => mm_interconnect_0_onchip_ram_s1_clken,                           --                                                                  .clken
			onchip_ram_s2_address                                                   => mm_interconnect_0_onchip_ram_s2_address,                         --                                                     onchip_ram_s2.address
			onchip_ram_s2_write                                                     => mm_interconnect_0_onchip_ram_s2_write,                           --                                                                  .write
			onchip_ram_s2_readdata                                                  => mm_interconnect_0_onchip_ram_s2_readdata,                        --                                                                  .readdata
			onchip_ram_s2_writedata                                                 => mm_interconnect_0_onchip_ram_s2_writedata,                       --                                                                  .writedata
			onchip_ram_s2_byteenable                                                => mm_interconnect_0_onchip_ram_s2_byteenable,                      --                                                                  .byteenable
			onchip_ram_s2_chipselect                                                => mm_interconnect_0_onchip_ram_s2_chipselect,                      --                                                                  .chipselect
			onchip_ram_s2_clken                                                     => mm_interconnect_0_onchip_ram_s2_clken,                           --                                                                  .clken
			pb_cpu_to_io_s0_address                                                 => mm_interconnect_0_pb_cpu_to_io_s0_address,                       --                                                   pb_cpu_to_io_s0.address
			pb_cpu_to_io_s0_write                                                   => mm_interconnect_0_pb_cpu_to_io_s0_write,                         --                                                                  .write
			pb_cpu_to_io_s0_read                                                    => mm_interconnect_0_pb_cpu_to_io_s0_read,                          --                                                                  .read
			pb_cpu_to_io_s0_readdata                                                => mm_interconnect_0_pb_cpu_to_io_s0_readdata,                      --                                                                  .readdata
			pb_cpu_to_io_s0_writedata                                               => mm_interconnect_0_pb_cpu_to_io_s0_writedata,                     --                                                                  .writedata
			pb_cpu_to_io_s0_burstcount                                              => mm_interconnect_0_pb_cpu_to_io_s0_burstcount,                    --                                                                  .burstcount
			pb_cpu_to_io_s0_byteenable                                              => mm_interconnect_0_pb_cpu_to_io_s0_byteenable,                    --                                                                  .byteenable
			pb_cpu_to_io_s0_readdatavalid                                           => mm_interconnect_0_pb_cpu_to_io_s0_readdatavalid,                 --                                                                  .readdatavalid
			pb_cpu_to_io_s0_waitrequest                                             => mm_interconnect_0_pb_cpu_to_io_s0_waitrequest,                   --                                                                  .waitrequest
			pb_cpu_to_io_s0_debugaccess                                             => mm_interconnect_0_pb_cpu_to_io_s0_debugaccess,                   --                                                                  .debugaccess
			sgdma_rx_csr_address                                                    => mm_interconnect_0_sgdma_rx_csr_address,                          --                                                      sgdma_rx_csr.address
			sgdma_rx_csr_write                                                      => mm_interconnect_0_sgdma_rx_csr_write,                            --                                                                  .write
			sgdma_rx_csr_read                                                       => mm_interconnect_0_sgdma_rx_csr_read,                             --                                                                  .read
			sgdma_rx_csr_readdata                                                   => mm_interconnect_0_sgdma_rx_csr_readdata,                         --                                                                  .readdata
			sgdma_rx_csr_writedata                                                  => mm_interconnect_0_sgdma_rx_csr_writedata,                        --                                                                  .writedata
			sgdma_rx_csr_chipselect                                                 => mm_interconnect_0_sgdma_rx_csr_chipselect,                       --                                                                  .chipselect
			sgdma_tx_csr_address                                                    => mm_interconnect_0_sgdma_tx_csr_address,                          --                                                      sgdma_tx_csr.address
			sgdma_tx_csr_write                                                      => mm_interconnect_0_sgdma_tx_csr_write,                            --                                                                  .write
			sgdma_tx_csr_read                                                       => mm_interconnect_0_sgdma_tx_csr_read,                             --                                                                  .read
			sgdma_tx_csr_readdata                                                   => mm_interconnect_0_sgdma_tx_csr_readdata,                         --                                                                  .readdata
			sgdma_tx_csr_writedata                                                  => mm_interconnect_0_sgdma_tx_csr_writedata,                        --                                                                  .writedata
			sgdma_tx_csr_chipselect                                                 => mm_interconnect_0_sgdma_tx_csr_chipselect,                       --                                                                  .chipselect
			tse_mac_control_port_address                                            => mm_interconnect_0_tse_mac_control_port_address,                  --                                              tse_mac_control_port.address
			tse_mac_control_port_write                                              => mm_interconnect_0_tse_mac_control_port_write,                    --                                                                  .write
			tse_mac_control_port_read                                               => mm_interconnect_0_tse_mac_control_port_read,                     --                                                                  .read
			tse_mac_control_port_readdata                                           => mm_interconnect_0_tse_mac_control_port_readdata,                 --                                                                  .readdata
			tse_mac_control_port_writedata                                          => mm_interconnect_0_tse_mac_control_port_writedata,                --                                                                  .writedata
			tse_mac_control_port_waitrequest                                        => mm_interconnect_0_tse_mac_control_port_waitrequest               --                                                                  .waitrequest
		);

	mm_interconnect_1 : component Nios_CPU_qsys_mm_interconnect_1
		port map (
			clkin_50_clk_clk                               => clk_clk,                                                     --                             clkin_50_clk.clk
			jtag_uart_0_reset_reset_bridge_in_reset_reset  => rst_controller_001_reset_out_reset,                          --  jtag_uart_0_reset_reset_bridge_in_reset.reset
			pb_cpu_to_io_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                              -- pb_cpu_to_io_reset_reset_bridge_in_reset.reset
			pb_cpu_to_io_m0_address                        => pb_cpu_to_io_m0_address,                                     --                          pb_cpu_to_io_m0.address
			pb_cpu_to_io_m0_waitrequest                    => pb_cpu_to_io_m0_waitrequest,                                 --                                         .waitrequest
			pb_cpu_to_io_m0_burstcount                     => pb_cpu_to_io_m0_burstcount,                                  --                                         .burstcount
			pb_cpu_to_io_m0_byteenable                     => pb_cpu_to_io_m0_byteenable,                                  --                                         .byteenable
			pb_cpu_to_io_m0_read                           => pb_cpu_to_io_m0_read,                                        --                                         .read
			pb_cpu_to_io_m0_readdata                       => pb_cpu_to_io_m0_readdata,                                    --                                         .readdata
			pb_cpu_to_io_m0_readdatavalid                  => pb_cpu_to_io_m0_readdatavalid,                               --                                         .readdatavalid
			pb_cpu_to_io_m0_write                          => pb_cpu_to_io_m0_write,                                       --                                         .write
			pb_cpu_to_io_m0_writedata                      => pb_cpu_to_io_m0_writedata,                                   --                                         .writedata
			pb_cpu_to_io_m0_debugaccess                    => pb_cpu_to_io_m0_debugaccess,                                 --                                         .debugaccess
			high_res_timer_s1_address                      => mm_interconnect_1_high_res_timer_s1_address,                 --                        high_res_timer_s1.address
			high_res_timer_s1_write                        => mm_interconnect_1_high_res_timer_s1_write,                   --                                         .write
			high_res_timer_s1_readdata                     => mm_interconnect_1_high_res_timer_s1_readdata,                --                                         .readdata
			high_res_timer_s1_writedata                    => mm_interconnect_1_high_res_timer_s1_writedata,               --                                         .writedata
			high_res_timer_s1_chipselect                   => mm_interconnect_1_high_res_timer_s1_chipselect,              --                                         .chipselect
			jtag_uart_0_avalon_jtag_slave_address          => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address,     --            jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write            => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write,       --                                         .write
			jtag_uart_0_avalon_jtag_slave_read             => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read,        --                                         .read
			jtag_uart_0_avalon_jtag_slave_readdata         => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata,    --                                         .readdata
			jtag_uart_0_avalon_jtag_slave_writedata        => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata,   --                                         .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest      => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest, --                                         .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect       => mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect,  --                                         .chipselect
			sys_clk_timer_s1_address                       => mm_interconnect_1_sys_clk_timer_s1_address,                  --                         sys_clk_timer_s1.address
			sys_clk_timer_s1_write                         => mm_interconnect_1_sys_clk_timer_s1_write,                    --                                         .write
			sys_clk_timer_s1_readdata                      => mm_interconnect_1_sys_clk_timer_s1_readdata,                 --                                         .readdata
			sys_clk_timer_s1_writedata                     => mm_interconnect_1_sys_clk_timer_s1_writedata,                --                                         .writedata
			sys_clk_timer_s1_chipselect                    => mm_interconnect_1_sys_clk_timer_s1_chipselect,               --                                         .chipselect
			sysid_control_slave_address                    => mm_interconnect_1_sysid_control_slave_address,               --                      sysid_control_slave.address
			sysid_control_slave_readdata                   => mm_interconnect_1_sysid_control_slave_readdata               --                                         .readdata
		);

	irq_mapper : component Nios_CPU_qsys_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,       -- receiver4.irq
			sender_irq    => cpu_irq_irq                     --    sender.irq
		);

	avalon_st_adapter : component Nios_CPU_qsys_avalon_st_adapter
		generic map (
			inBitsPerSymbol => 8,
			inUsePackets    => 1,
			inDataWidth     => 32,
			inChannelWidth  => 0,
			inErrorWidth    => 6,
			inUseEmptyPort  => 1,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 2,
			outDataWidth    => 32,
			outChannelWidth => 0,
			outErrorWidth   => 6,
			outUseEmptyPort => 1,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk        => clk_clk,                               -- in_clk_0.clk
			in_rst_0_reset      => rst_controller_001_reset_out_reset,    -- in_rst_0.reset
			in_0_data           => tse_mac_receive_data,                  --     in_0.data
			in_0_valid          => tse_mac_receive_valid,                 --         .valid
			in_0_ready          => tse_mac_receive_ready,                 --         .ready
			in_0_startofpacket  => tse_mac_receive_startofpacket,         --         .startofpacket
			in_0_endofpacket    => tse_mac_receive_endofpacket,           --         .endofpacket
			in_0_empty          => tse_mac_receive_empty,                 --         .empty
			in_0_error          => tse_mac_receive_error,                 --         .error
			out_0_data          => avalon_st_adapter_out_0_data,          --    out_0.data
			out_0_valid         => avalon_st_adapter_out_0_valid,         --         .valid
			out_0_ready         => avalon_st_adapter_out_0_ready,         --         .ready
			out_0_startofpacket => avalon_st_adapter_out_0_startofpacket, --         .startofpacket
			out_0_endofpacket   => avalon_st_adapter_out_0_endofpacket,   --         .endofpacket
			out_0_empty         => avalon_st_adapter_out_0_empty,         --         .empty
			out_0_error         => avalon_st_adapter_out_0_error          --         .error
		);

	rst_controller : component nios_cpu_qsys_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 3,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => merged_resets_in_reset_reset_n_ports_inv, -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,            -- reset_in1.reset
			reset_in2      => merged_resets_in_reset_reset_n_ports_inv, -- reset_in2.reset
			clk            => clk_clk,                                  --       clk.clk
			reset_out      => rst_controller_reset_out_reset,           -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,       --          .reset_req
			reset_req_in0  => '0',                                      -- (terminated)
			reset_req_in1  => '0',                                      -- (terminated)
			reset_req_in2  => '0',                                      -- (terminated)
			reset_in3      => '0',                                      -- (terminated)
			reset_req_in3  => '0',                                      -- (terminated)
			reset_in4      => '0',                                      -- (terminated)
			reset_req_in4  => '0',                                      -- (terminated)
			reset_in5      => '0',                                      -- (terminated)
			reset_req_in5  => '0',                                      -- (terminated)
			reset_in6      => '0',                                      -- (terminated)
			reset_req_in6  => '0',                                      -- (terminated)
			reset_in7      => '0',                                      -- (terminated)
			reset_req_in7  => '0',                                      -- (terminated)
			reset_in8      => '0',                                      -- (terminated)
			reset_req_in8  => '0',                                      -- (terminated)
			reset_in9      => '0',                                      -- (terminated)
			reset_req_in9  => '0',                                      -- (terminated)
			reset_in10     => '0',                                      -- (terminated)
			reset_req_in10 => '0',                                      -- (terminated)
			reset_in11     => '0',                                      -- (terminated)
			reset_req_in11 => '0',                                      -- (terminated)
			reset_in12     => '0',                                      -- (terminated)
			reset_req_in12 => '0',                                      -- (terminated)
			reset_in13     => '0',                                      -- (terminated)
			reset_req_in13 => '0',                                      -- (terminated)
			reset_in14     => '0',                                      -- (terminated)
			reset_req_in14 => '0',                                      -- (terminated)
			reset_in15     => '0',                                      -- (terminated)
			reset_req_in15 => '0'                                       -- (terminated)
		);

	rst_controller_001 : component nios_cpu_qsys_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => merged_resets_in_reset_reset_n_ports_inv, -- reset_in0.reset
			reset_in1      => merged_resets_in_reset_reset_n_ports_inv, -- reset_in1.reset
			clk            => clk_clk,                                  --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,       -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req,   --          .reset_req
			reset_req_in0  => '0',                                      -- (terminated)
			reset_req_in1  => '0',                                      -- (terminated)
			reset_in2      => '0',                                      -- (terminated)
			reset_req_in2  => '0',                                      -- (terminated)
			reset_in3      => '0',                                      -- (terminated)
			reset_req_in3  => '0',                                      -- (terminated)
			reset_in4      => '0',                                      -- (terminated)
			reset_req_in4  => '0',                                      -- (terminated)
			reset_in5      => '0',                                      -- (terminated)
			reset_req_in5  => '0',                                      -- (terminated)
			reset_in6      => '0',                                      -- (terminated)
			reset_req_in6  => '0',                                      -- (terminated)
			reset_in7      => '0',                                      -- (terminated)
			reset_req_in7  => '0',                                      -- (terminated)
			reset_in8      => '0',                                      -- (terminated)
			reset_req_in8  => '0',                                      -- (terminated)
			reset_in9      => '0',                                      -- (terminated)
			reset_req_in9  => '0',                                      -- (terminated)
			reset_in10     => '0',                                      -- (terminated)
			reset_req_in10 => '0',                                      -- (terminated)
			reset_in11     => '0',                                      -- (terminated)
			reset_req_in11 => '0',                                      -- (terminated)
			reset_in12     => '0',                                      -- (terminated)
			reset_req_in12 => '0',                                      -- (terminated)
			reset_in13     => '0',                                      -- (terminated)
			reset_req_in13 => '0',                                      -- (terminated)
			reset_in14     => '0',                                      -- (terminated)
			reset_req_in14 => '0',                                      -- (terminated)
			reset_in15     => '0',                                      -- (terminated)
			reset_req_in15 => '0'                                       -- (terminated)
		);

	rst_controller_002 : component nios_cpu_qsys_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => merged_resets_in_reset_reset_n_ports_inv, -- reset_in0.reset
			clk            => mem_if_lpddr2_emif_0_afi_clk_clk,         --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,       -- reset_out.reset
			reset_req      => open,                                     -- (terminated)
			reset_req_in0  => '0',                                      -- (terminated)
			reset_in1      => '0',                                      -- (terminated)
			reset_req_in1  => '0',                                      -- (terminated)
			reset_in2      => '0',                                      -- (terminated)
			reset_req_in2  => '0',                                      -- (terminated)
			reset_in3      => '0',                                      -- (terminated)
			reset_req_in3  => '0',                                      -- (terminated)
			reset_in4      => '0',                                      -- (terminated)
			reset_req_in4  => '0',                                      -- (terminated)
			reset_in5      => '0',                                      -- (terminated)
			reset_req_in5  => '0',                                      -- (terminated)
			reset_in6      => '0',                                      -- (terminated)
			reset_req_in6  => '0',                                      -- (terminated)
			reset_in7      => '0',                                      -- (terminated)
			reset_req_in7  => '0',                                      -- (terminated)
			reset_in8      => '0',                                      -- (terminated)
			reset_req_in8  => '0',                                      -- (terminated)
			reset_in9      => '0',                                      -- (terminated)
			reset_req_in9  => '0',                                      -- (terminated)
			reset_in10     => '0',                                      -- (terminated)
			reset_req_in10 => '0',                                      -- (terminated)
			reset_in11     => '0',                                      -- (terminated)
			reset_req_in11 => '0',                                      -- (terminated)
			reset_in12     => '0',                                      -- (terminated)
			reset_req_in12 => '0',                                      -- (terminated)
			reset_in13     => '0',                                      -- (terminated)
			reset_req_in13 => '0',                                      -- (terminated)
			reset_in14     => '0',                                      -- (terminated)
			reset_req_in14 => '0',                                      -- (terminated)
			reset_in15     => '0',                                      -- (terminated)
			reset_req_in15 => '0'                                       -- (terminated)
		);

	merged_resets_in_reset_reset_n_ports_inv <= not merged_resets_in_reset_reset_n;

	mm_interconnect_0_mem_if_lpddr2_emif_0_avl_0_inv <= not mem_if_lpddr2_emif_0_avl_0_waitrequest;

	mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_1_sys_clk_timer_s1_write_ports_inv <= not mm_interconnect_1_sys_clk_timer_s1_write;

	mm_interconnect_1_high_res_timer_s1_write_ports_inv <= not mm_interconnect_1_high_res_timer_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of Nios_CPU_qsys
