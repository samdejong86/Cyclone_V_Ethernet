// Nios_CPU_qsys.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module Nios_CPU_qsys (
		output wire [26:0] cfi_flash_atb_bridge_0_out_tcm_address_out,      //          cfi_flash_atb_bridge_0_out.tcm_address_out
		output wire [0:0]  cfi_flash_atb_bridge_0_out_tcm_read_n_out,       //                                    .tcm_read_n_out
		output wire [0:0]  cfi_flash_atb_bridge_0_out_tcm_write_n_out,      //                                    .tcm_write_n_out
		inout  wire [15:0] cfi_flash_atb_bridge_0_out_tcm_data_out,         //                                    .tcm_data_out
		output wire [0:0]  cfi_flash_atb_bridge_0_out_tcm_chipselect_n_out, //                                    .tcm_chipselect_n_out
		input  wire        clk_clk,                                         //                                 clk.clk
		input  wire        merged_resets_in_reset_reset_n,                  //              merged_resets_in_reset.reset_n
		input  wire [7:0]  tse_mac_mac_gmii_connection_gmii_rx_d,           //         tse_mac_mac_gmii_connection.gmii_rx_d
		input  wire        tse_mac_mac_gmii_connection_gmii_rx_dv,          //                                    .gmii_rx_dv
		input  wire        tse_mac_mac_gmii_connection_gmii_rx_err,         //                                    .gmii_rx_err
		output wire [7:0]  tse_mac_mac_gmii_connection_gmii_tx_d,           //                                    .gmii_tx_d
		output wire        tse_mac_mac_gmii_connection_gmii_tx_en,          //                                    .gmii_tx_en
		output wire        tse_mac_mac_gmii_connection_gmii_tx_err,         //                                    .gmii_tx_err
		output wire        tse_mac_mac_mdio_connection_mdc,                 //         tse_mac_mac_mdio_connection.mdc
		input  wire        tse_mac_mac_mdio_connection_mdio_in,             //                                    .mdio_in
		output wire        tse_mac_mac_mdio_connection_mdio_out,            //                                    .mdio_out
		output wire        tse_mac_mac_mdio_connection_mdio_oen,            //                                    .mdio_oen
		input  wire [3:0]  tse_mac_mac_mii_connection_mii_rx_d,             //          tse_mac_mac_mii_connection.mii_rx_d
		input  wire        tse_mac_mac_mii_connection_mii_rx_dv,            //                                    .mii_rx_dv
		input  wire        tse_mac_mac_mii_connection_mii_rx_err,           //                                    .mii_rx_err
		output wire [3:0]  tse_mac_mac_mii_connection_mii_tx_d,             //                                    .mii_tx_d
		output wire        tse_mac_mac_mii_connection_mii_tx_en,            //                                    .mii_tx_en
		output wire        tse_mac_mac_mii_connection_mii_tx_err,           //                                    .mii_tx_err
		input  wire        tse_mac_mac_mii_connection_mii_crs,              //                                    .mii_crs
		input  wire        tse_mac_mac_mii_connection_mii_col,              //                                    .mii_col
		input  wire        tse_mac_mac_misc_connection_xon_gen,             //         tse_mac_mac_misc_connection.xon_gen
		input  wire        tse_mac_mac_misc_connection_xoff_gen,            //                                    .xoff_gen
		input  wire        tse_mac_mac_misc_connection_ff_tx_crc_fwd,       //                                    .ff_tx_crc_fwd
		output wire        tse_mac_mac_misc_connection_ff_tx_septy,         //                                    .ff_tx_septy
		output wire        tse_mac_mac_misc_connection_tx_ff_uflow,         //                                    .tx_ff_uflow
		output wire        tse_mac_mac_misc_connection_ff_tx_a_full,        //                                    .ff_tx_a_full
		output wire        tse_mac_mac_misc_connection_ff_tx_a_empty,       //                                    .ff_tx_a_empty
		output wire [17:0] tse_mac_mac_misc_connection_rx_err_stat,         //                                    .rx_err_stat
		output wire [3:0]  tse_mac_mac_misc_connection_rx_frm_type,         //                                    .rx_frm_type
		output wire        tse_mac_mac_misc_connection_ff_rx_dsav,          //                                    .ff_rx_dsav
		output wire        tse_mac_mac_misc_connection_ff_rx_a_full,        //                                    .ff_rx_a_full
		output wire        tse_mac_mac_misc_connection_ff_rx_a_empty,       //                                    .ff_rx_a_empty
		input  wire        tse_mac_mac_status_connection_set_10,            //       tse_mac_mac_status_connection.set_10
		input  wire        tse_mac_mac_status_connection_set_1000,          //                                    .set_1000
		output wire        tse_mac_mac_status_connection_eth_mode,          //                                    .eth_mode
		output wire        tse_mac_mac_status_connection_ena_10,            //                                    .ena_10
		input  wire        tse_mac_pcs_mac_rx_clock_connection_clk,         // tse_mac_pcs_mac_rx_clock_connection.clk
		input  wire        tse_mac_pcs_mac_tx_clock_connection_clk          // tse_mac_pcs_mac_tx_clock_connection.clk
	);

	wire         sgdma_tx_out_valid;                                          // sgdma_tx:out_valid -> tse_mac:ff_tx_wren
	wire  [31:0] sgdma_tx_out_data;                                           // sgdma_tx:out_data -> tse_mac:ff_tx_data
	wire         sgdma_tx_out_ready;                                          // tse_mac:ff_tx_rdy -> sgdma_tx:out_ready
	wire         sgdma_tx_out_startofpacket;                                  // sgdma_tx:out_startofpacket -> tse_mac:ff_tx_sop
	wire         sgdma_tx_out_endofpacket;                                    // sgdma_tx:out_endofpacket -> tse_mac:ff_tx_eop
	wire         sgdma_tx_out_error;                                          // sgdma_tx:out_error -> tse_mac:ff_tx_err
	wire   [1:0] sgdma_tx_out_empty;                                          // sgdma_tx:out_empty -> tse_mac:ff_tx_mod
	wire         ext_flash_tcm_data_outen;                                    // ext_flash:tcm_data_outen -> cfi_flash_atb_bridge_0:tcs_tcm_data_outen
	wire         ext_flash_tcm_request;                                       // ext_flash:tcm_request -> cfi_flash_atb_bridge_0:request
	wire         ext_flash_tcm_write_n_out;                                   // ext_flash:tcm_write_n_out -> cfi_flash_atb_bridge_0:tcs_tcm_write_n_out
	wire         ext_flash_tcm_read_n_out;                                    // ext_flash:tcm_read_n_out -> cfi_flash_atb_bridge_0:tcs_tcm_read_n_out
	wire         ext_flash_tcm_grant;                                         // cfi_flash_atb_bridge_0:grant -> ext_flash:tcm_grant
	wire         ext_flash_tcm_chipselect_n_out;                              // ext_flash:tcm_chipselect_n_out -> cfi_flash_atb_bridge_0:tcs_tcm_chipselect_n_out
	wire  [26:0] ext_flash_tcm_address_out;                                   // ext_flash:tcm_address_out -> cfi_flash_atb_bridge_0:tcs_tcm_address_out
	wire  [15:0] ext_flash_tcm_data_out;                                      // ext_flash:tcm_data_out -> cfi_flash_atb_bridge_0:tcs_tcm_data_out
	wire  [15:0] ext_flash_tcm_data_in;                                       // cfi_flash_atb_bridge_0:tcs_tcm_data_in -> ext_flash:tcm_data_in
	wire  [31:0] cpu_data_master_readdata;                                    // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                 // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                 // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [27:0] cpu_data_master_address;                                     // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                  // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                        // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_readdatavalid;                               // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire         cpu_data_master_write;                                       // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                   // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                             // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                          // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [27:0] cpu_instruction_master_address;                              // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                 // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                        // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire  [31:0] sgdma_tx_m_read_readdata;                                    // mm_interconnect_0:sgdma_tx_m_read_readdata -> sgdma_tx:m_read_readdata
	wire         sgdma_tx_m_read_waitrequest;                                 // mm_interconnect_0:sgdma_tx_m_read_waitrequest -> sgdma_tx:m_read_waitrequest
	wire  [31:0] sgdma_tx_m_read_address;                                     // sgdma_tx:m_read_address -> mm_interconnect_0:sgdma_tx_m_read_address
	wire         sgdma_tx_m_read_read;                                        // sgdma_tx:m_read_read -> mm_interconnect_0:sgdma_tx_m_read_read
	wire         sgdma_tx_m_read_readdatavalid;                               // mm_interconnect_0:sgdma_tx_m_read_readdatavalid -> sgdma_tx:m_read_readdatavalid
	wire         sgdma_rx_m_write_waitrequest;                                // mm_interconnect_0:sgdma_rx_m_write_waitrequest -> sgdma_rx:m_write_waitrequest
	wire  [31:0] sgdma_rx_m_write_address;                                    // sgdma_rx:m_write_address -> mm_interconnect_0:sgdma_rx_m_write_address
	wire   [3:0] sgdma_rx_m_write_byteenable;                                 // sgdma_rx:m_write_byteenable -> mm_interconnect_0:sgdma_rx_m_write_byteenable
	wire         sgdma_rx_m_write_write;                                      // sgdma_rx:m_write_write -> mm_interconnect_0:sgdma_rx_m_write_write
	wire  [31:0] sgdma_rx_m_write_writedata;                                  // sgdma_rx:m_write_writedata -> mm_interconnect_0:sgdma_rx_m_write_writedata
	wire  [31:0] sgdma_rx_descriptor_read_readdata;                           // mm_interconnect_0:sgdma_rx_descriptor_read_readdata -> sgdma_rx:descriptor_read_readdata
	wire         sgdma_rx_descriptor_read_waitrequest;                        // mm_interconnect_0:sgdma_rx_descriptor_read_waitrequest -> sgdma_rx:descriptor_read_waitrequest
	wire  [31:0] sgdma_rx_descriptor_read_address;                            // sgdma_rx:descriptor_read_address -> mm_interconnect_0:sgdma_rx_descriptor_read_address
	wire         sgdma_rx_descriptor_read_read;                               // sgdma_rx:descriptor_read_read -> mm_interconnect_0:sgdma_rx_descriptor_read_read
	wire         sgdma_rx_descriptor_read_readdatavalid;                      // mm_interconnect_0:sgdma_rx_descriptor_read_readdatavalid -> sgdma_rx:descriptor_read_readdatavalid
	wire  [31:0] sgdma_tx_descriptor_read_readdata;                           // mm_interconnect_0:sgdma_tx_descriptor_read_readdata -> sgdma_tx:descriptor_read_readdata
	wire         sgdma_tx_descriptor_read_waitrequest;                        // mm_interconnect_0:sgdma_tx_descriptor_read_waitrequest -> sgdma_tx:descriptor_read_waitrequest
	wire  [31:0] sgdma_tx_descriptor_read_address;                            // sgdma_tx:descriptor_read_address -> mm_interconnect_0:sgdma_tx_descriptor_read_address
	wire         sgdma_tx_descriptor_read_read;                               // sgdma_tx:descriptor_read_read -> mm_interconnect_0:sgdma_tx_descriptor_read_read
	wire         sgdma_tx_descriptor_read_readdatavalid;                      // mm_interconnect_0:sgdma_tx_descriptor_read_readdatavalid -> sgdma_tx:descriptor_read_readdatavalid
	wire         sgdma_rx_descriptor_write_waitrequest;                       // mm_interconnect_0:sgdma_rx_descriptor_write_waitrequest -> sgdma_rx:descriptor_write_waitrequest
	wire  [31:0] sgdma_rx_descriptor_write_address;                           // sgdma_rx:descriptor_write_address -> mm_interconnect_0:sgdma_rx_descriptor_write_address
	wire         sgdma_rx_descriptor_write_write;                             // sgdma_rx:descriptor_write_write -> mm_interconnect_0:sgdma_rx_descriptor_write_write
	wire  [31:0] sgdma_rx_descriptor_write_writedata;                         // sgdma_rx:descriptor_write_writedata -> mm_interconnect_0:sgdma_rx_descriptor_write_writedata
	wire         sgdma_tx_descriptor_write_waitrequest;                       // mm_interconnect_0:sgdma_tx_descriptor_write_waitrequest -> sgdma_tx:descriptor_write_waitrequest
	wire  [31:0] sgdma_tx_descriptor_write_address;                           // sgdma_tx:descriptor_write_address -> mm_interconnect_0:sgdma_tx_descriptor_write_address
	wire         sgdma_tx_descriptor_write_write;                             // sgdma_tx:descriptor_write_write -> mm_interconnect_0:sgdma_tx_descriptor_write_write
	wire  [31:0] sgdma_tx_descriptor_write_writedata;                         // sgdma_tx:descriptor_write_writedata -> mm_interconnect_0:sgdma_tx_descriptor_write_writedata
	wire  [31:0] mm_interconnect_0_tse_mac_control_port_readdata;             // tse_mac:reg_data_out -> mm_interconnect_0:tse_mac_control_port_readdata
	wire         mm_interconnect_0_tse_mac_control_port_waitrequest;          // tse_mac:reg_busy -> mm_interconnect_0:tse_mac_control_port_waitrequest
	wire   [7:0] mm_interconnect_0_tse_mac_control_port_address;              // mm_interconnect_0:tse_mac_control_port_address -> tse_mac:reg_addr
	wire         mm_interconnect_0_tse_mac_control_port_read;                 // mm_interconnect_0:tse_mac_control_port_read -> tse_mac:reg_rd
	wire         mm_interconnect_0_tse_mac_control_port_write;                // mm_interconnect_0:tse_mac_control_port_write -> tse_mac:reg_wr
	wire  [31:0] mm_interconnect_0_tse_mac_control_port_writedata;            // mm_interconnect_0:tse_mac_control_port_writedata -> tse_mac:reg_data_in
	wire         mm_interconnect_0_sgdma_tx_csr_chipselect;                   // mm_interconnect_0:sgdma_tx_csr_chipselect -> sgdma_tx:csr_chipselect
	wire  [31:0] mm_interconnect_0_sgdma_tx_csr_readdata;                     // sgdma_tx:csr_readdata -> mm_interconnect_0:sgdma_tx_csr_readdata
	wire   [3:0] mm_interconnect_0_sgdma_tx_csr_address;                      // mm_interconnect_0:sgdma_tx_csr_address -> sgdma_tx:csr_address
	wire         mm_interconnect_0_sgdma_tx_csr_read;                         // mm_interconnect_0:sgdma_tx_csr_read -> sgdma_tx:csr_read
	wire         mm_interconnect_0_sgdma_tx_csr_write;                        // mm_interconnect_0:sgdma_tx_csr_write -> sgdma_tx:csr_write
	wire  [31:0] mm_interconnect_0_sgdma_tx_csr_writedata;                    // mm_interconnect_0:sgdma_tx_csr_writedata -> sgdma_tx:csr_writedata
	wire         mm_interconnect_0_sgdma_rx_csr_chipselect;                   // mm_interconnect_0:sgdma_rx_csr_chipselect -> sgdma_rx:csr_chipselect
	wire  [31:0] mm_interconnect_0_sgdma_rx_csr_readdata;                     // sgdma_rx:csr_readdata -> mm_interconnect_0:sgdma_rx_csr_readdata
	wire   [3:0] mm_interconnect_0_sgdma_rx_csr_address;                      // mm_interconnect_0:sgdma_rx_csr_address -> sgdma_rx:csr_address
	wire         mm_interconnect_0_sgdma_rx_csr_read;                         // mm_interconnect_0:sgdma_rx_csr_read -> sgdma_rx:csr_read
	wire         mm_interconnect_0_sgdma_rx_csr_write;                        // mm_interconnect_0:sgdma_rx_csr_write -> sgdma_rx:csr_write
	wire  [31:0] mm_interconnect_0_sgdma_rx_csr_writedata;                    // mm_interconnect_0:sgdma_rx_csr_writedata -> sgdma_rx:csr_writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;              // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;           // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;           // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;               // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                  // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;            // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;                 // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;             // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_pb_cpu_to_io_s0_readdata;                  // pb_cpu_to_io:s0_readdata -> mm_interconnect_0:pb_cpu_to_io_s0_readdata
	wire         mm_interconnect_0_pb_cpu_to_io_s0_waitrequest;               // pb_cpu_to_io:s0_waitrequest -> mm_interconnect_0:pb_cpu_to_io_s0_waitrequest
	wire         mm_interconnect_0_pb_cpu_to_io_s0_debugaccess;               // mm_interconnect_0:pb_cpu_to_io_s0_debugaccess -> pb_cpu_to_io:s0_debugaccess
	wire   [9:0] mm_interconnect_0_pb_cpu_to_io_s0_address;                   // mm_interconnect_0:pb_cpu_to_io_s0_address -> pb_cpu_to_io:s0_address
	wire         mm_interconnect_0_pb_cpu_to_io_s0_read;                      // mm_interconnect_0:pb_cpu_to_io_s0_read -> pb_cpu_to_io:s0_read
	wire   [3:0] mm_interconnect_0_pb_cpu_to_io_s0_byteenable;                // mm_interconnect_0:pb_cpu_to_io_s0_byteenable -> pb_cpu_to_io:s0_byteenable
	wire         mm_interconnect_0_pb_cpu_to_io_s0_readdatavalid;             // pb_cpu_to_io:s0_readdatavalid -> mm_interconnect_0:pb_cpu_to_io_s0_readdatavalid
	wire         mm_interconnect_0_pb_cpu_to_io_s0_write;                     // mm_interconnect_0:pb_cpu_to_io_s0_write -> pb_cpu_to_io:s0_write
	wire  [31:0] mm_interconnect_0_pb_cpu_to_io_s0_writedata;                 // mm_interconnect_0:pb_cpu_to_io_s0_writedata -> pb_cpu_to_io:s0_writedata
	wire   [0:0] mm_interconnect_0_pb_cpu_to_io_s0_burstcount;                // mm_interconnect_0:pb_cpu_to_io_s0_burstcount -> pb_cpu_to_io:s0_burstcount
	wire         mm_interconnect_0_onchip_ram_s1_chipselect;                  // mm_interconnect_0:onchip_ram_s1_chipselect -> onchip_ram:chipselect
	wire  [31:0] mm_interconnect_0_onchip_ram_s1_readdata;                    // onchip_ram:readdata -> mm_interconnect_0:onchip_ram_s1_readdata
	wire  [18:0] mm_interconnect_0_onchip_ram_s1_address;                     // mm_interconnect_0:onchip_ram_s1_address -> onchip_ram:address
	wire   [3:0] mm_interconnect_0_onchip_ram_s1_byteenable;                  // mm_interconnect_0:onchip_ram_s1_byteenable -> onchip_ram:byteenable
	wire         mm_interconnect_0_onchip_ram_s1_write;                       // mm_interconnect_0:onchip_ram_s1_write -> onchip_ram:write
	wire  [31:0] mm_interconnect_0_onchip_ram_s1_writedata;                   // mm_interconnect_0:onchip_ram_s1_writedata -> onchip_ram:writedata
	wire         mm_interconnect_0_onchip_ram_s1_clken;                       // mm_interconnect_0:onchip_ram_s1_clken -> onchip_ram:clken
	wire         mm_interconnect_0_descriptor_memory_s1_chipselect;           // mm_interconnect_0:descriptor_memory_s1_chipselect -> descriptor_memory:chipselect
	wire  [31:0] mm_interconnect_0_descriptor_memory_s1_readdata;             // descriptor_memory:readdata -> mm_interconnect_0:descriptor_memory_s1_readdata
	wire  [10:0] mm_interconnect_0_descriptor_memory_s1_address;              // mm_interconnect_0:descriptor_memory_s1_address -> descriptor_memory:address
	wire   [3:0] mm_interconnect_0_descriptor_memory_s1_byteenable;           // mm_interconnect_0:descriptor_memory_s1_byteenable -> descriptor_memory:byteenable
	wire         mm_interconnect_0_descriptor_memory_s1_write;                // mm_interconnect_0:descriptor_memory_s1_write -> descriptor_memory:write
	wire  [31:0] mm_interconnect_0_descriptor_memory_s1_writedata;            // mm_interconnect_0:descriptor_memory_s1_writedata -> descriptor_memory:writedata
	wire         mm_interconnect_0_descriptor_memory_s1_clken;                // mm_interconnect_0:descriptor_memory_s1_clken -> descriptor_memory:clken
	wire         mm_interconnect_0_onchip_ram_s2_chipselect;                  // mm_interconnect_0:onchip_ram_s2_chipselect -> onchip_ram:chipselect2
	wire  [31:0] mm_interconnect_0_onchip_ram_s2_readdata;                    // onchip_ram:readdata2 -> mm_interconnect_0:onchip_ram_s2_readdata
	wire  [18:0] mm_interconnect_0_onchip_ram_s2_address;                     // mm_interconnect_0:onchip_ram_s2_address -> onchip_ram:address2
	wire   [3:0] mm_interconnect_0_onchip_ram_s2_byteenable;                  // mm_interconnect_0:onchip_ram_s2_byteenable -> onchip_ram:byteenable2
	wire         mm_interconnect_0_onchip_ram_s2_write;                       // mm_interconnect_0:onchip_ram_s2_write -> onchip_ram:write2
	wire  [31:0] mm_interconnect_0_onchip_ram_s2_writedata;                   // mm_interconnect_0:onchip_ram_s2_writedata -> onchip_ram:writedata2
	wire         mm_interconnect_0_onchip_ram_s2_clken;                       // mm_interconnect_0:onchip_ram_s2_clken -> onchip_ram:clken2
	wire  [15:0] mm_interconnect_0_ext_flash_uas_readdata;                    // ext_flash:uas_readdata -> mm_interconnect_0:ext_flash_uas_readdata
	wire         mm_interconnect_0_ext_flash_uas_waitrequest;                 // ext_flash:uas_waitrequest -> mm_interconnect_0:ext_flash_uas_waitrequest
	wire         mm_interconnect_0_ext_flash_uas_debugaccess;                 // mm_interconnect_0:ext_flash_uas_debugaccess -> ext_flash:uas_debugaccess
	wire  [26:0] mm_interconnect_0_ext_flash_uas_address;                     // mm_interconnect_0:ext_flash_uas_address -> ext_flash:uas_address
	wire         mm_interconnect_0_ext_flash_uas_read;                        // mm_interconnect_0:ext_flash_uas_read -> ext_flash:uas_read
	wire   [1:0] mm_interconnect_0_ext_flash_uas_byteenable;                  // mm_interconnect_0:ext_flash_uas_byteenable -> ext_flash:uas_byteenable
	wire         mm_interconnect_0_ext_flash_uas_readdatavalid;               // ext_flash:uas_readdatavalid -> mm_interconnect_0:ext_flash_uas_readdatavalid
	wire         mm_interconnect_0_ext_flash_uas_lock;                        // mm_interconnect_0:ext_flash_uas_lock -> ext_flash:uas_lock
	wire         mm_interconnect_0_ext_flash_uas_write;                       // mm_interconnect_0:ext_flash_uas_write -> ext_flash:uas_write
	wire  [15:0] mm_interconnect_0_ext_flash_uas_writedata;                   // mm_interconnect_0:ext_flash_uas_writedata -> ext_flash:uas_writedata
	wire   [1:0] mm_interconnect_0_ext_flash_uas_burstcount;                  // mm_interconnect_0:ext_flash_uas_burstcount -> ext_flash:uas_burstcount
	wire         pb_cpu_to_io_m0_waitrequest;                                 // mm_interconnect_1:pb_cpu_to_io_m0_waitrequest -> pb_cpu_to_io:m0_waitrequest
	wire  [31:0] pb_cpu_to_io_m0_readdata;                                    // mm_interconnect_1:pb_cpu_to_io_m0_readdata -> pb_cpu_to_io:m0_readdata
	wire         pb_cpu_to_io_m0_debugaccess;                                 // pb_cpu_to_io:m0_debugaccess -> mm_interconnect_1:pb_cpu_to_io_m0_debugaccess
	wire   [9:0] pb_cpu_to_io_m0_address;                                     // pb_cpu_to_io:m0_address -> mm_interconnect_1:pb_cpu_to_io_m0_address
	wire         pb_cpu_to_io_m0_read;                                        // pb_cpu_to_io:m0_read -> mm_interconnect_1:pb_cpu_to_io_m0_read
	wire   [3:0] pb_cpu_to_io_m0_byteenable;                                  // pb_cpu_to_io:m0_byteenable -> mm_interconnect_1:pb_cpu_to_io_m0_byteenable
	wire         pb_cpu_to_io_m0_readdatavalid;                               // mm_interconnect_1:pb_cpu_to_io_m0_readdatavalid -> pb_cpu_to_io:m0_readdatavalid
	wire  [31:0] pb_cpu_to_io_m0_writedata;                                   // pb_cpu_to_io:m0_writedata -> mm_interconnect_1:pb_cpu_to_io_m0_writedata
	wire         pb_cpu_to_io_m0_write;                                       // pb_cpu_to_io:m0_write -> mm_interconnect_1:pb_cpu_to_io_m0_write
	wire   [0:0] pb_cpu_to_io_m0_burstcount;                                  // pb_cpu_to_io:m0_burstcount -> mm_interconnect_1:pb_cpu_to_io_m0_burstcount
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_1:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;              // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;               // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire         mm_interconnect_1_sys_clk_timer_s1_chipselect;               // mm_interconnect_1:sys_clk_timer_s1_chipselect -> sys_clk_timer:chipselect
	wire  [15:0] mm_interconnect_1_sys_clk_timer_s1_readdata;                 // sys_clk_timer:readdata -> mm_interconnect_1:sys_clk_timer_s1_readdata
	wire   [2:0] mm_interconnect_1_sys_clk_timer_s1_address;                  // mm_interconnect_1:sys_clk_timer_s1_address -> sys_clk_timer:address
	wire         mm_interconnect_1_sys_clk_timer_s1_write;                    // mm_interconnect_1:sys_clk_timer_s1_write -> sys_clk_timer:write_n
	wire  [15:0] mm_interconnect_1_sys_clk_timer_s1_writedata;                // mm_interconnect_1:sys_clk_timer_s1_writedata -> sys_clk_timer:writedata
	wire         mm_interconnect_1_high_res_timer_s1_chipselect;              // mm_interconnect_1:high_res_timer_s1_chipselect -> high_res_timer:chipselect
	wire  [15:0] mm_interconnect_1_high_res_timer_s1_readdata;                // high_res_timer:readdata -> mm_interconnect_1:high_res_timer_s1_readdata
	wire   [2:0] mm_interconnect_1_high_res_timer_s1_address;                 // mm_interconnect_1:high_res_timer_s1_address -> high_res_timer:address
	wire         mm_interconnect_1_high_res_timer_s1_write;                   // mm_interconnect_1:high_res_timer_s1_write -> high_res_timer:write_n
	wire  [15:0] mm_interconnect_1_high_res_timer_s1_writedata;               // mm_interconnect_1:high_res_timer_s1_writedata -> high_res_timer:writedata
	wire         irq_mapper_receiver0_irq;                                    // sgdma_rx:csr_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // sgdma_tx:csr_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // sys_clk_timer:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                    // high_res_timer:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver4_irq
	wire  [31:0] cpu_irq_irq;                                                 // irq_mapper:sender_irq -> cpu:irq
	wire         tse_mac_receive_valid;                                       // tse_mac:ff_rx_dval -> avalon_st_adapter:in_0_valid
	wire  [31:0] tse_mac_receive_data;                                        // tse_mac:ff_rx_data -> avalon_st_adapter:in_0_data
	wire         tse_mac_receive_ready;                                       // avalon_st_adapter:in_0_ready -> tse_mac:ff_rx_rdy
	wire         tse_mac_receive_startofpacket;                               // tse_mac:ff_rx_sop -> avalon_st_adapter:in_0_startofpacket
	wire         tse_mac_receive_endofpacket;                                 // tse_mac:ff_rx_eop -> avalon_st_adapter:in_0_endofpacket
	wire   [5:0] tse_mac_receive_error;                                       // tse_mac:rx_err -> avalon_st_adapter:in_0_error
	wire   [1:0] tse_mac_receive_empty;                                       // tse_mac:ff_rx_mod -> avalon_st_adapter:in_0_empty
	wire         avalon_st_adapter_out_0_valid;                               // avalon_st_adapter:out_0_valid -> sgdma_rx:in_valid
	wire  [31:0] avalon_st_adapter_out_0_data;                                // avalon_st_adapter:out_0_data -> sgdma_rx:in_data
	wire         avalon_st_adapter_out_0_ready;                               // sgdma_rx:in_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                       // avalon_st_adapter:out_0_startofpacket -> sgdma_rx:in_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                         // avalon_st_adapter:out_0_endofpacket -> sgdma_rx:in_endofpacket
	wire   [5:0] avalon_st_adapter_out_0_error;                               // avalon_st_adapter:out_0_error -> sgdma_rx:in_error
	wire   [1:0] avalon_st_adapter_out_0_empty;                               // avalon_st_adapter:out_0_empty -> sgdma_rx:in_empty
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, cfi_flash_atb_bridge_0:reset, descriptor_memory:reset, ext_flash:reset_reset, high_res_timer:reset_n, jtag_uart_0:rst_n, mm_interconnect_0:sgdma_tx_reset_reset_bridge_in_reset_reset, mm_interconnect_1:jtag_uart_0_reset_reset_bridge_in_reset_reset, onchip_ram:reset, onchip_ram:reset2, rst_translator:in_reset, sgdma_rx:system_reset_n, sgdma_tx:system_reset_n, sys_clk_timer:reset_n, sysid:reset_n, tse_mac:reset]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [descriptor_memory:reset_req, onchip_ram:reset_req, onchip_ram:reset_req2, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [cpu:reset_n, irq_mapper:reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, mm_interconnect_1:pb_cpu_to_io_reset_reset_bridge_in_reset_reset, pb_cpu_to_io:reset, rst_translator_001:in_reset]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [cpu:reset_req, rst_translator_001:reset_req_in]
	wire         cpu_debug_reset_request_reset;                               // cpu:debug_reset_request -> rst_controller_001:reset_in1

	Nios_CPU_qsys_cfi_flash_atb_bridge_0 cfi_flash_atb_bridge_0 (
		.clk                      (clk_clk),                                         //   clk.clk
		.reset                    (rst_controller_reset_out_reset),                  // reset.reset
		.request                  (ext_flash_tcm_request),                           //   tcs.request
		.grant                    (ext_flash_tcm_grant),                             //      .grant
		.tcs_tcm_address_out      (ext_flash_tcm_address_out),                       //      .address_out
		.tcs_tcm_read_n_out       (ext_flash_tcm_read_n_out),                        //      .read_n_out
		.tcs_tcm_write_n_out      (ext_flash_tcm_write_n_out),                       //      .write_n_out
		.tcs_tcm_data_out         (ext_flash_tcm_data_out),                          //      .data_out
		.tcs_tcm_data_outen       (ext_flash_tcm_data_outen),                        //      .data_outen
		.tcs_tcm_data_in          (ext_flash_tcm_data_in),                           //      .data_in
		.tcs_tcm_chipselect_n_out (ext_flash_tcm_chipselect_n_out),                  //      .chipselect_n_out
		.tcm_address_out          (cfi_flash_atb_bridge_0_out_tcm_address_out),      //   out.tcm_address_out
		.tcm_read_n_out           (cfi_flash_atb_bridge_0_out_tcm_read_n_out),       //      .tcm_read_n_out
		.tcm_write_n_out          (cfi_flash_atb_bridge_0_out_tcm_write_n_out),      //      .tcm_write_n_out
		.tcm_data_out             (cfi_flash_atb_bridge_0_out_tcm_data_out),         //      .tcm_data_out
		.tcm_chipselect_n_out     (cfi_flash_atb_bridge_0_out_tcm_chipselect_n_out)  //      .tcm_chipselect_n_out
	);

	Nios_CPU_qsys_cpu cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),               //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),            //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	Nios_CPU_qsys_descriptor_memory descriptor_memory (
		.clk        (clk_clk),                                           //   clk1.clk
		.address    (mm_interconnect_0_descriptor_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_descriptor_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_descriptor_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_descriptor_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_descriptor_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_descriptor_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_descriptor_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                    // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),                //       .reset_req
		.freeze     (1'b0)                                               // (terminated)
	);

	Nios_CPU_qsys_ext_flash #(
		.TCM_ADDRESS_W                  (27),
		.TCM_DATA_W                     (16),
		.TCM_BYTEENABLE_W               (2),
		.TCM_READ_WAIT                  (135),
		.TCM_WRITE_WAIT                 (135),
		.TCM_SETUP_WAIT                 (25),
		.TCM_DATA_HOLD                  (20),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (2),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (0),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (0),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (1)
	) ext_flash (
		.clk_clk              (clk_clk),                                       //   clk.clk
		.reset_reset          (rst_controller_reset_out_reset),                // reset.reset
		.uas_address          (mm_interconnect_0_ext_flash_uas_address),       //   uas.address
		.uas_burstcount       (mm_interconnect_0_ext_flash_uas_burstcount),    //      .burstcount
		.uas_read             (mm_interconnect_0_ext_flash_uas_read),          //      .read
		.uas_write            (mm_interconnect_0_ext_flash_uas_write),         //      .write
		.uas_waitrequest      (mm_interconnect_0_ext_flash_uas_waitrequest),   //      .waitrequest
		.uas_readdatavalid    (mm_interconnect_0_ext_flash_uas_readdatavalid), //      .readdatavalid
		.uas_byteenable       (mm_interconnect_0_ext_flash_uas_byteenable),    //      .byteenable
		.uas_readdata         (mm_interconnect_0_ext_flash_uas_readdata),      //      .readdata
		.uas_writedata        (mm_interconnect_0_ext_flash_uas_writedata),     //      .writedata
		.uas_lock             (mm_interconnect_0_ext_flash_uas_lock),          //      .lock
		.uas_debugaccess      (mm_interconnect_0_ext_flash_uas_debugaccess),   //      .debugaccess
		.tcm_write_n_out      (ext_flash_tcm_write_n_out),                     //   tcm.write_n_out
		.tcm_read_n_out       (ext_flash_tcm_read_n_out),                      //      .read_n_out
		.tcm_chipselect_n_out (ext_flash_tcm_chipselect_n_out),                //      .chipselect_n_out
		.tcm_request          (ext_flash_tcm_request),                         //      .request
		.tcm_grant            (ext_flash_tcm_grant),                           //      .grant
		.tcm_address_out      (ext_flash_tcm_address_out),                     //      .address_out
		.tcm_data_out         (ext_flash_tcm_data_out),                        //      .data_out
		.tcm_data_outen       (ext_flash_tcm_data_outen),                      //      .data_outen
		.tcm_data_in          (ext_flash_tcm_data_in)                          //      .data_in
	);

	Nios_CPU_qsys_high_res_timer high_res_timer (
		.clk        (clk_clk),                                        //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                // reset.reset_n
		.address    (mm_interconnect_1_high_res_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_high_res_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_high_res_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_high_res_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_high_res_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                        //   irq.irq
	);

	Nios_CPU_qsys_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver4_irq)                                     //               irq.irq
	);

	Nios_CPU_qsys_onchip_ram onchip_ram (
		.clk         (clk_clk),                                    //   clk1.clk
		.address     (mm_interconnect_0_onchip_ram_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_onchip_ram_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_onchip_ram_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_onchip_ram_s1_write),      //       .write
		.readdata    (mm_interconnect_0_onchip_ram_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_onchip_ram_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_onchip_ram_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),         //       .reset_req
		.address2    (mm_interconnect_0_onchip_ram_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_onchip_ram_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_onchip_ram_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_onchip_ram_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_onchip_ram_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_onchip_ram_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_onchip_ram_s2_byteenable), //       .byteenable
		.clk2        (clk_clk),                                    //   clk2.clk
		.reset2      (rst_controller_reset_out_reset),             // reset2.reset
		.reset_req2  (rst_controller_reset_out_reset_req),         //       .reset_req
		.freeze      (1'b0)                                        // (terminated)
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (10),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) pb_cpu_to_io (
		.clk              (clk_clk),                                         //   clk.clk
		.reset            (rst_controller_001_reset_out_reset),              // reset.reset
		.s0_waitrequest   (mm_interconnect_0_pb_cpu_to_io_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_pb_cpu_to_io_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_pb_cpu_to_io_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_pb_cpu_to_io_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_pb_cpu_to_io_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_pb_cpu_to_io_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_pb_cpu_to_io_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_pb_cpu_to_io_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_pb_cpu_to_io_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_pb_cpu_to_io_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (pb_cpu_to_io_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (pb_cpu_to_io_m0_readdata),                        //      .readdata
		.m0_readdatavalid (pb_cpu_to_io_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (pb_cpu_to_io_m0_burstcount),                      //      .burstcount
		.m0_writedata     (pb_cpu_to_io_m0_writedata),                       //      .writedata
		.m0_address       (pb_cpu_to_io_m0_address),                         //      .address
		.m0_write         (pb_cpu_to_io_m0_write),                           //      .write
		.m0_read          (pb_cpu_to_io_m0_read),                            //      .read
		.m0_byteenable    (pb_cpu_to_io_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (pb_cpu_to_io_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                                // (terminated)
		.m0_response      (2'b00)                                            // (terminated)
	);

	Nios_CPU_qsys_sgdma_rx sgdma_rx (
		.clk                           (clk_clk),                                   //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),           //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_sgdma_rx_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_sgdma_rx_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_sgdma_rx_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_sgdma_rx_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_sgdma_rx_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_sgdma_rx_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_rx_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_rx_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_rx_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (sgdma_rx_descriptor_read_address),          //                 .address
		.descriptor_read_read          (sgdma_rx_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (sgdma_rx_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_rx_descriptor_write_address),         //                 .address
		.descriptor_write_write        (sgdma_rx_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (sgdma_rx_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver0_irq),                  //          csr_irq.irq
		.in_startofpacket              (avalon_st_adapter_out_0_startofpacket),     //               in.startofpacket
		.in_endofpacket                (avalon_st_adapter_out_0_endofpacket),       //                 .endofpacket
		.in_data                       (avalon_st_adapter_out_0_data),              //                 .data
		.in_valid                      (avalon_st_adapter_out_0_valid),             //                 .valid
		.in_ready                      (avalon_st_adapter_out_0_ready),             //                 .ready
		.in_empty                      (avalon_st_adapter_out_0_empty),             //                 .empty
		.in_error                      (avalon_st_adapter_out_0_error),             //                 .error
		.m_write_waitrequest           (sgdma_rx_m_write_waitrequest),              //          m_write.waitrequest
		.m_write_address               (sgdma_rx_m_write_address),                  //                 .address
		.m_write_write                 (sgdma_rx_m_write_write),                    //                 .write
		.m_write_writedata             (sgdma_rx_m_write_writedata),                //                 .writedata
		.m_write_byteenable            (sgdma_rx_m_write_byteenable)                //                 .byteenable
	);

	Nios_CPU_qsys_sgdma_tx sgdma_tx (
		.clk                           (clk_clk),                                   //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),           //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_sgdma_tx_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_sgdma_tx_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_sgdma_tx_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_sgdma_tx_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_sgdma_tx_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_sgdma_tx_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (sgdma_tx_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (sgdma_tx_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (sgdma_tx_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (sgdma_tx_descriptor_read_address),          //                 .address
		.descriptor_read_read          (sgdma_tx_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (sgdma_tx_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (sgdma_tx_descriptor_write_address),         //                 .address
		.descriptor_write_write        (sgdma_tx_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (sgdma_tx_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver1_irq),                  //          csr_irq.irq
		.m_read_readdata               (sgdma_tx_m_read_readdata),                  //           m_read.readdata
		.m_read_readdatavalid          (sgdma_tx_m_read_readdatavalid),             //                 .readdatavalid
		.m_read_waitrequest            (sgdma_tx_m_read_waitrequest),               //                 .waitrequest
		.m_read_address                (sgdma_tx_m_read_address),                   //                 .address
		.m_read_read                   (sgdma_tx_m_read_read),                      //                 .read
		.out_data                      (sgdma_tx_out_data),                         //              out.data
		.out_valid                     (sgdma_tx_out_valid),                        //                 .valid
		.out_ready                     (sgdma_tx_out_ready),                        //                 .ready
		.out_endofpacket               (sgdma_tx_out_endofpacket),                  //                 .endofpacket
		.out_startofpacket             (sgdma_tx_out_startofpacket),                //                 .startofpacket
		.out_empty                     (sgdma_tx_out_empty),                        //                 .empty
		.out_error                     (sgdma_tx_out_error)                         //                 .error
	);

	Nios_CPU_qsys_sys_clk_timer sys_clk_timer (
		.clk        (clk_clk),                                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               // reset.reset_n
		.address    (mm_interconnect_1_sys_clk_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_sys_clk_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_sys_clk_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_sys_clk_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_sys_clk_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                       //   irq.irq
	);

	Nios_CPU_qsys_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	Nios_CPU_qsys_tse_mac tse_mac (
		.clk           (clk_clk),                                            // control_port_clock_connection.clk
		.reset         (rst_controller_reset_out_reset),                     //              reset_connection.reset
		.reg_addr      (mm_interconnect_0_tse_mac_control_port_address),     //                  control_port.address
		.reg_data_out  (mm_interconnect_0_tse_mac_control_port_readdata),    //                              .readdata
		.reg_rd        (mm_interconnect_0_tse_mac_control_port_read),        //                              .read
		.reg_data_in   (mm_interconnect_0_tse_mac_control_port_writedata),   //                              .writedata
		.reg_wr        (mm_interconnect_0_tse_mac_control_port_write),       //                              .write
		.reg_busy      (mm_interconnect_0_tse_mac_control_port_waitrequest), //                              .waitrequest
		.tx_clk        (tse_mac_pcs_mac_tx_clock_connection_clk),            //   pcs_mac_tx_clock_connection.clk
		.rx_clk        (tse_mac_pcs_mac_rx_clock_connection_clk),            //   pcs_mac_rx_clock_connection.clk
		.set_10        (tse_mac_mac_status_connection_set_10),               //         mac_status_connection.set_10
		.set_1000      (tse_mac_mac_status_connection_set_1000),             //                              .set_1000
		.eth_mode      (tse_mac_mac_status_connection_eth_mode),             //                              .eth_mode
		.ena_10        (tse_mac_mac_status_connection_ena_10),               //                              .ena_10
		.gm_rx_d       (tse_mac_mac_gmii_connection_gmii_rx_d),              //           mac_gmii_connection.gmii_rx_d
		.gm_rx_dv      (tse_mac_mac_gmii_connection_gmii_rx_dv),             //                              .gmii_rx_dv
		.gm_rx_err     (tse_mac_mac_gmii_connection_gmii_rx_err),            //                              .gmii_rx_err
		.gm_tx_d       (tse_mac_mac_gmii_connection_gmii_tx_d),              //                              .gmii_tx_d
		.gm_tx_en      (tse_mac_mac_gmii_connection_gmii_tx_en),             //                              .gmii_tx_en
		.gm_tx_err     (tse_mac_mac_gmii_connection_gmii_tx_err),            //                              .gmii_tx_err
		.m_rx_d        (tse_mac_mac_mii_connection_mii_rx_d),                //            mac_mii_connection.mii_rx_d
		.m_rx_en       (tse_mac_mac_mii_connection_mii_rx_dv),               //                              .mii_rx_dv
		.m_rx_err      (tse_mac_mac_mii_connection_mii_rx_err),              //                              .mii_rx_err
		.m_tx_d        (tse_mac_mac_mii_connection_mii_tx_d),                //                              .mii_tx_d
		.m_tx_en       (tse_mac_mac_mii_connection_mii_tx_en),               //                              .mii_tx_en
		.m_tx_err      (tse_mac_mac_mii_connection_mii_tx_err),              //                              .mii_tx_err
		.m_rx_crs      (tse_mac_mac_mii_connection_mii_crs),                 //                              .mii_crs
		.m_rx_col      (tse_mac_mac_mii_connection_mii_col),                 //                              .mii_col
		.ff_rx_clk     (clk_clk),                                            //      receive_clock_connection.clk
		.ff_tx_clk     (clk_clk),                                            //     transmit_clock_connection.clk
		.ff_rx_data    (tse_mac_receive_data),                               //                       receive.data
		.ff_rx_eop     (tse_mac_receive_endofpacket),                        //                              .endofpacket
		.rx_err        (tse_mac_receive_error),                              //                              .error
		.ff_rx_mod     (tse_mac_receive_empty),                              //                              .empty
		.ff_rx_rdy     (tse_mac_receive_ready),                              //                              .ready
		.ff_rx_sop     (tse_mac_receive_startofpacket),                      //                              .startofpacket
		.ff_rx_dval    (tse_mac_receive_valid),                              //                              .valid
		.ff_tx_data    (sgdma_tx_out_data),                                  //                      transmit.data
		.ff_tx_eop     (sgdma_tx_out_endofpacket),                           //                              .endofpacket
		.ff_tx_err     (sgdma_tx_out_error),                                 //                              .error
		.ff_tx_mod     (sgdma_tx_out_empty),                                 //                              .empty
		.ff_tx_rdy     (sgdma_tx_out_ready),                                 //                              .ready
		.ff_tx_sop     (sgdma_tx_out_startofpacket),                         //                              .startofpacket
		.ff_tx_wren    (sgdma_tx_out_valid),                                 //                              .valid
		.mdc           (tse_mac_mac_mdio_connection_mdc),                    //           mac_mdio_connection.mdc
		.mdio_in       (tse_mac_mac_mdio_connection_mdio_in),                //                              .mdio_in
		.mdio_out      (tse_mac_mac_mdio_connection_mdio_out),               //                              .mdio_out
		.mdio_oen      (tse_mac_mac_mdio_connection_mdio_oen),               //                              .mdio_oen
		.xon_gen       (tse_mac_mac_misc_connection_xon_gen),                //           mac_misc_connection.xon_gen
		.xoff_gen      (tse_mac_mac_misc_connection_xoff_gen),               //                              .xoff_gen
		.ff_tx_crc_fwd (tse_mac_mac_misc_connection_ff_tx_crc_fwd),          //                              .ff_tx_crc_fwd
		.ff_tx_septy   (tse_mac_mac_misc_connection_ff_tx_septy),            //                              .ff_tx_septy
		.tx_ff_uflow   (tse_mac_mac_misc_connection_tx_ff_uflow),            //                              .tx_ff_uflow
		.ff_tx_a_full  (tse_mac_mac_misc_connection_ff_tx_a_full),           //                              .ff_tx_a_full
		.ff_tx_a_empty (tse_mac_mac_misc_connection_ff_tx_a_empty),          //                              .ff_tx_a_empty
		.rx_err_stat   (tse_mac_mac_misc_connection_rx_err_stat),            //                              .rx_err_stat
		.rx_frm_type   (tse_mac_mac_misc_connection_rx_frm_type),            //                              .rx_frm_type
		.ff_rx_dsav    (tse_mac_mac_misc_connection_ff_rx_dsav),             //                              .ff_rx_dsav
		.ff_rx_a_full  (tse_mac_mac_misc_connection_ff_rx_a_full),           //                              .ff_rx_a_full
		.ff_rx_a_empty (tse_mac_mac_misc_connection_ff_rx_a_empty)           //                              .ff_rx_a_empty
	);

	Nios_CPU_qsys_mm_interconnect_0 mm_interconnect_0 (
		.clkin_50_clk_clk                           (clk_clk),                                            //                         clkin_50_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset      (rst_controller_001_reset_out_reset),                 //      cpu_reset_reset_bridge_in_reset.reset
		.sgdma_tx_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                     // sgdma_tx_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                    (cpu_data_master_address),                            //                      cpu_data_master.address
		.cpu_data_master_waitrequest                (cpu_data_master_waitrequest),                        //                                     .waitrequest
		.cpu_data_master_byteenable                 (cpu_data_master_byteenable),                         //                                     .byteenable
		.cpu_data_master_read                       (cpu_data_master_read),                               //                                     .read
		.cpu_data_master_readdata                   (cpu_data_master_readdata),                           //                                     .readdata
		.cpu_data_master_readdatavalid              (cpu_data_master_readdatavalid),                      //                                     .readdatavalid
		.cpu_data_master_write                      (cpu_data_master_write),                              //                                     .write
		.cpu_data_master_writedata                  (cpu_data_master_writedata),                          //                                     .writedata
		.cpu_data_master_debugaccess                (cpu_data_master_debugaccess),                        //                                     .debugaccess
		.cpu_instruction_master_address             (cpu_instruction_master_address),                     //               cpu_instruction_master.address
		.cpu_instruction_master_waitrequest         (cpu_instruction_master_waitrequest),                 //                                     .waitrequest
		.cpu_instruction_master_read                (cpu_instruction_master_read),                        //                                     .read
		.cpu_instruction_master_readdata            (cpu_instruction_master_readdata),                    //                                     .readdata
		.cpu_instruction_master_readdatavalid       (cpu_instruction_master_readdatavalid),               //                                     .readdatavalid
		.sgdma_rx_descriptor_read_address           (sgdma_rx_descriptor_read_address),                   //             sgdma_rx_descriptor_read.address
		.sgdma_rx_descriptor_read_waitrequest       (sgdma_rx_descriptor_read_waitrequest),               //                                     .waitrequest
		.sgdma_rx_descriptor_read_read              (sgdma_rx_descriptor_read_read),                      //                                     .read
		.sgdma_rx_descriptor_read_readdata          (sgdma_rx_descriptor_read_readdata),                  //                                     .readdata
		.sgdma_rx_descriptor_read_readdatavalid     (sgdma_rx_descriptor_read_readdatavalid),             //                                     .readdatavalid
		.sgdma_rx_descriptor_write_address          (sgdma_rx_descriptor_write_address),                  //            sgdma_rx_descriptor_write.address
		.sgdma_rx_descriptor_write_waitrequest      (sgdma_rx_descriptor_write_waitrequest),              //                                     .waitrequest
		.sgdma_rx_descriptor_write_write            (sgdma_rx_descriptor_write_write),                    //                                     .write
		.sgdma_rx_descriptor_write_writedata        (sgdma_rx_descriptor_write_writedata),                //                                     .writedata
		.sgdma_rx_m_write_address                   (sgdma_rx_m_write_address),                           //                     sgdma_rx_m_write.address
		.sgdma_rx_m_write_waitrequest               (sgdma_rx_m_write_waitrequest),                       //                                     .waitrequest
		.sgdma_rx_m_write_byteenable                (sgdma_rx_m_write_byteenable),                        //                                     .byteenable
		.sgdma_rx_m_write_write                     (sgdma_rx_m_write_write),                             //                                     .write
		.sgdma_rx_m_write_writedata                 (sgdma_rx_m_write_writedata),                         //                                     .writedata
		.sgdma_tx_descriptor_read_address           (sgdma_tx_descriptor_read_address),                   //             sgdma_tx_descriptor_read.address
		.sgdma_tx_descriptor_read_waitrequest       (sgdma_tx_descriptor_read_waitrequest),               //                                     .waitrequest
		.sgdma_tx_descriptor_read_read              (sgdma_tx_descriptor_read_read),                      //                                     .read
		.sgdma_tx_descriptor_read_readdata          (sgdma_tx_descriptor_read_readdata),                  //                                     .readdata
		.sgdma_tx_descriptor_read_readdatavalid     (sgdma_tx_descriptor_read_readdatavalid),             //                                     .readdatavalid
		.sgdma_tx_descriptor_write_address          (sgdma_tx_descriptor_write_address),                  //            sgdma_tx_descriptor_write.address
		.sgdma_tx_descriptor_write_waitrequest      (sgdma_tx_descriptor_write_waitrequest),              //                                     .waitrequest
		.sgdma_tx_descriptor_write_write            (sgdma_tx_descriptor_write_write),                    //                                     .write
		.sgdma_tx_descriptor_write_writedata        (sgdma_tx_descriptor_write_writedata),                //                                     .writedata
		.sgdma_tx_m_read_address                    (sgdma_tx_m_read_address),                            //                      sgdma_tx_m_read.address
		.sgdma_tx_m_read_waitrequest                (sgdma_tx_m_read_waitrequest),                        //                                     .waitrequest
		.sgdma_tx_m_read_read                       (sgdma_tx_m_read_read),                               //                                     .read
		.sgdma_tx_m_read_readdata                   (sgdma_tx_m_read_readdata),                           //                                     .readdata
		.sgdma_tx_m_read_readdatavalid              (sgdma_tx_m_read_readdatavalid),                      //                                     .readdatavalid
		.cpu_debug_mem_slave_address                (mm_interconnect_0_cpu_debug_mem_slave_address),      //                  cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                  (mm_interconnect_0_cpu_debug_mem_slave_write),        //                                     .write
		.cpu_debug_mem_slave_read                   (mm_interconnect_0_cpu_debug_mem_slave_read),         //                                     .read
		.cpu_debug_mem_slave_readdata               (mm_interconnect_0_cpu_debug_mem_slave_readdata),     //                                     .readdata
		.cpu_debug_mem_slave_writedata              (mm_interconnect_0_cpu_debug_mem_slave_writedata),    //                                     .writedata
		.cpu_debug_mem_slave_byteenable             (mm_interconnect_0_cpu_debug_mem_slave_byteenable),   //                                     .byteenable
		.cpu_debug_mem_slave_waitrequest            (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),  //                                     .waitrequest
		.cpu_debug_mem_slave_debugaccess            (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),  //                                     .debugaccess
		.descriptor_memory_s1_address               (mm_interconnect_0_descriptor_memory_s1_address),     //                 descriptor_memory_s1.address
		.descriptor_memory_s1_write                 (mm_interconnect_0_descriptor_memory_s1_write),       //                                     .write
		.descriptor_memory_s1_readdata              (mm_interconnect_0_descriptor_memory_s1_readdata),    //                                     .readdata
		.descriptor_memory_s1_writedata             (mm_interconnect_0_descriptor_memory_s1_writedata),   //                                     .writedata
		.descriptor_memory_s1_byteenable            (mm_interconnect_0_descriptor_memory_s1_byteenable),  //                                     .byteenable
		.descriptor_memory_s1_chipselect            (mm_interconnect_0_descriptor_memory_s1_chipselect),  //                                     .chipselect
		.descriptor_memory_s1_clken                 (mm_interconnect_0_descriptor_memory_s1_clken),       //                                     .clken
		.ext_flash_uas_address                      (mm_interconnect_0_ext_flash_uas_address),            //                        ext_flash_uas.address
		.ext_flash_uas_write                        (mm_interconnect_0_ext_flash_uas_write),              //                                     .write
		.ext_flash_uas_read                         (mm_interconnect_0_ext_flash_uas_read),               //                                     .read
		.ext_flash_uas_readdata                     (mm_interconnect_0_ext_flash_uas_readdata),           //                                     .readdata
		.ext_flash_uas_writedata                    (mm_interconnect_0_ext_flash_uas_writedata),          //                                     .writedata
		.ext_flash_uas_burstcount                   (mm_interconnect_0_ext_flash_uas_burstcount),         //                                     .burstcount
		.ext_flash_uas_byteenable                   (mm_interconnect_0_ext_flash_uas_byteenable),         //                                     .byteenable
		.ext_flash_uas_readdatavalid                (mm_interconnect_0_ext_flash_uas_readdatavalid),      //                                     .readdatavalid
		.ext_flash_uas_waitrequest                  (mm_interconnect_0_ext_flash_uas_waitrequest),        //                                     .waitrequest
		.ext_flash_uas_lock                         (mm_interconnect_0_ext_flash_uas_lock),               //                                     .lock
		.ext_flash_uas_debugaccess                  (mm_interconnect_0_ext_flash_uas_debugaccess),        //                                     .debugaccess
		.onchip_ram_s1_address                      (mm_interconnect_0_onchip_ram_s1_address),            //                        onchip_ram_s1.address
		.onchip_ram_s1_write                        (mm_interconnect_0_onchip_ram_s1_write),              //                                     .write
		.onchip_ram_s1_readdata                     (mm_interconnect_0_onchip_ram_s1_readdata),           //                                     .readdata
		.onchip_ram_s1_writedata                    (mm_interconnect_0_onchip_ram_s1_writedata),          //                                     .writedata
		.onchip_ram_s1_byteenable                   (mm_interconnect_0_onchip_ram_s1_byteenable),         //                                     .byteenable
		.onchip_ram_s1_chipselect                   (mm_interconnect_0_onchip_ram_s1_chipselect),         //                                     .chipselect
		.onchip_ram_s1_clken                        (mm_interconnect_0_onchip_ram_s1_clken),              //                                     .clken
		.onchip_ram_s2_address                      (mm_interconnect_0_onchip_ram_s2_address),            //                        onchip_ram_s2.address
		.onchip_ram_s2_write                        (mm_interconnect_0_onchip_ram_s2_write),              //                                     .write
		.onchip_ram_s2_readdata                     (mm_interconnect_0_onchip_ram_s2_readdata),           //                                     .readdata
		.onchip_ram_s2_writedata                    (mm_interconnect_0_onchip_ram_s2_writedata),          //                                     .writedata
		.onchip_ram_s2_byteenable                   (mm_interconnect_0_onchip_ram_s2_byteenable),         //                                     .byteenable
		.onchip_ram_s2_chipselect                   (mm_interconnect_0_onchip_ram_s2_chipselect),         //                                     .chipselect
		.onchip_ram_s2_clken                        (mm_interconnect_0_onchip_ram_s2_clken),              //                                     .clken
		.pb_cpu_to_io_s0_address                    (mm_interconnect_0_pb_cpu_to_io_s0_address),          //                      pb_cpu_to_io_s0.address
		.pb_cpu_to_io_s0_write                      (mm_interconnect_0_pb_cpu_to_io_s0_write),            //                                     .write
		.pb_cpu_to_io_s0_read                       (mm_interconnect_0_pb_cpu_to_io_s0_read),             //                                     .read
		.pb_cpu_to_io_s0_readdata                   (mm_interconnect_0_pb_cpu_to_io_s0_readdata),         //                                     .readdata
		.pb_cpu_to_io_s0_writedata                  (mm_interconnect_0_pb_cpu_to_io_s0_writedata),        //                                     .writedata
		.pb_cpu_to_io_s0_burstcount                 (mm_interconnect_0_pb_cpu_to_io_s0_burstcount),       //                                     .burstcount
		.pb_cpu_to_io_s0_byteenable                 (mm_interconnect_0_pb_cpu_to_io_s0_byteenable),       //                                     .byteenable
		.pb_cpu_to_io_s0_readdatavalid              (mm_interconnect_0_pb_cpu_to_io_s0_readdatavalid),    //                                     .readdatavalid
		.pb_cpu_to_io_s0_waitrequest                (mm_interconnect_0_pb_cpu_to_io_s0_waitrequest),      //                                     .waitrequest
		.pb_cpu_to_io_s0_debugaccess                (mm_interconnect_0_pb_cpu_to_io_s0_debugaccess),      //                                     .debugaccess
		.sgdma_rx_csr_address                       (mm_interconnect_0_sgdma_rx_csr_address),             //                         sgdma_rx_csr.address
		.sgdma_rx_csr_write                         (mm_interconnect_0_sgdma_rx_csr_write),               //                                     .write
		.sgdma_rx_csr_read                          (mm_interconnect_0_sgdma_rx_csr_read),                //                                     .read
		.sgdma_rx_csr_readdata                      (mm_interconnect_0_sgdma_rx_csr_readdata),            //                                     .readdata
		.sgdma_rx_csr_writedata                     (mm_interconnect_0_sgdma_rx_csr_writedata),           //                                     .writedata
		.sgdma_rx_csr_chipselect                    (mm_interconnect_0_sgdma_rx_csr_chipselect),          //                                     .chipselect
		.sgdma_tx_csr_address                       (mm_interconnect_0_sgdma_tx_csr_address),             //                         sgdma_tx_csr.address
		.sgdma_tx_csr_write                         (mm_interconnect_0_sgdma_tx_csr_write),               //                                     .write
		.sgdma_tx_csr_read                          (mm_interconnect_0_sgdma_tx_csr_read),                //                                     .read
		.sgdma_tx_csr_readdata                      (mm_interconnect_0_sgdma_tx_csr_readdata),            //                                     .readdata
		.sgdma_tx_csr_writedata                     (mm_interconnect_0_sgdma_tx_csr_writedata),           //                                     .writedata
		.sgdma_tx_csr_chipselect                    (mm_interconnect_0_sgdma_tx_csr_chipselect),          //                                     .chipselect
		.tse_mac_control_port_address               (mm_interconnect_0_tse_mac_control_port_address),     //                 tse_mac_control_port.address
		.tse_mac_control_port_write                 (mm_interconnect_0_tse_mac_control_port_write),       //                                     .write
		.tse_mac_control_port_read                  (mm_interconnect_0_tse_mac_control_port_read),        //                                     .read
		.tse_mac_control_port_readdata              (mm_interconnect_0_tse_mac_control_port_readdata),    //                                     .readdata
		.tse_mac_control_port_writedata             (mm_interconnect_0_tse_mac_control_port_writedata),   //                                     .writedata
		.tse_mac_control_port_waitrequest           (mm_interconnect_0_tse_mac_control_port_waitrequest)  //                                     .waitrequest
	);

	Nios_CPU_qsys_mm_interconnect_1 mm_interconnect_1 (
		.clkin_50_clk_clk                               (clk_clk),                                                     //                             clkin_50_clk.clk
		.jtag_uart_0_reset_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),                              //  jtag_uart_0_reset_reset_bridge_in_reset.reset
		.pb_cpu_to_io_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // pb_cpu_to_io_reset_reset_bridge_in_reset.reset
		.pb_cpu_to_io_m0_address                        (pb_cpu_to_io_m0_address),                                     //                          pb_cpu_to_io_m0.address
		.pb_cpu_to_io_m0_waitrequest                    (pb_cpu_to_io_m0_waitrequest),                                 //                                         .waitrequest
		.pb_cpu_to_io_m0_burstcount                     (pb_cpu_to_io_m0_burstcount),                                  //                                         .burstcount
		.pb_cpu_to_io_m0_byteenable                     (pb_cpu_to_io_m0_byteenable),                                  //                                         .byteenable
		.pb_cpu_to_io_m0_read                           (pb_cpu_to_io_m0_read),                                        //                                         .read
		.pb_cpu_to_io_m0_readdata                       (pb_cpu_to_io_m0_readdata),                                    //                                         .readdata
		.pb_cpu_to_io_m0_readdatavalid                  (pb_cpu_to_io_m0_readdatavalid),                               //                                         .readdatavalid
		.pb_cpu_to_io_m0_write                          (pb_cpu_to_io_m0_write),                                       //                                         .write
		.pb_cpu_to_io_m0_writedata                      (pb_cpu_to_io_m0_writedata),                                   //                                         .writedata
		.pb_cpu_to_io_m0_debugaccess                    (pb_cpu_to_io_m0_debugaccess),                                 //                                         .debugaccess
		.high_res_timer_s1_address                      (mm_interconnect_1_high_res_timer_s1_address),                 //                        high_res_timer_s1.address
		.high_res_timer_s1_write                        (mm_interconnect_1_high_res_timer_s1_write),                   //                                         .write
		.high_res_timer_s1_readdata                     (mm_interconnect_1_high_res_timer_s1_readdata),                //                                         .readdata
		.high_res_timer_s1_writedata                    (mm_interconnect_1_high_res_timer_s1_writedata),               //                                         .writedata
		.high_res_timer_s1_chipselect                   (mm_interconnect_1_high_res_timer_s1_chipselect),              //                                         .chipselect
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_1_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.sys_clk_timer_s1_address                       (mm_interconnect_1_sys_clk_timer_s1_address),                  //                         sys_clk_timer_s1.address
		.sys_clk_timer_s1_write                         (mm_interconnect_1_sys_clk_timer_s1_write),                    //                                         .write
		.sys_clk_timer_s1_readdata                      (mm_interconnect_1_sys_clk_timer_s1_readdata),                 //                                         .readdata
		.sys_clk_timer_s1_writedata                     (mm_interconnect_1_sys_clk_timer_s1_writedata),                //                                         .writedata
		.sys_clk_timer_s1_chipselect                    (mm_interconnect_1_sys_clk_timer_s1_chipselect),               //                                         .chipselect
		.sysid_control_slave_address                    (mm_interconnect_1_sysid_control_slave_address),               //                      sysid_control_slave.address
		.sysid_control_slave_readdata                   (mm_interconnect_1_sysid_control_slave_readdata)               //                                         .readdata
	);

	Nios_CPU_qsys_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.sender_irq    (cpu_irq_irq)                         //    sender.irq
	);

	Nios_CPU_qsys_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (6),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (2),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (6),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (clk_clk),                               // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),        // in_rst_0.reset
		.in_0_data           (tse_mac_receive_data),                  //     in_0.data
		.in_0_valid          (tse_mac_receive_valid),                 //         .valid
		.in_0_ready          (tse_mac_receive_ready),                 //         .ready
		.in_0_startofpacket  (tse_mac_receive_startofpacket),         //         .startofpacket
		.in_0_endofpacket    (tse_mac_receive_endofpacket),           //         .endofpacket
		.in_0_empty          (tse_mac_receive_empty),                 //         .empty
		.in_0_error          (tse_mac_receive_error),                 //         .error
		.out_0_data          (avalon_st_adapter_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty),         //         .empty
		.out_0_error         (avalon_st_adapter_out_0_error)          //         .error
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~merged_resets_in_reset_reset_n),    // reset_in0.reset
		.reset_in1      (~merged_resets_in_reset_reset_n),    // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (3),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~merged_resets_in_reset_reset_n),        // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),          // reset_in1.reset
		.reset_in2      (~merged_resets_in_reset_reset_n),        // reset_in2.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
