-- eth_std_main_system.vhd

-- Generated using ACDS version 16.1 196

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity eth_std_main_system is
	port (
		button_pio_external_connection_export       : in    std_logic_vector(2 downto 0)  := (others => '0'); -- button_pio_external_connection.export
		clk_125_clk_in_clk                          : in    std_logic                     := '0';             --                 clk_125_clk_in.clk
		clk_125_clk_in_reset_reset_n                : in    std_logic                     := '0';             --           clk_125_clk_in_reset.reset_n
		clk_50_clk_in_clk                           : in    std_logic                     := '0';             --                  clk_50_clk_in.clk
		clk_50_clk_in_reset_reset_n                 : in    std_logic                     := '0';             --            clk_50_clk_in_reset.reset_n
		ddr2_top_memory_mem_ca                      : out   std_logic_vector(9 downto 0);                     --                ddr2_top_memory.mem_ca
		ddr2_top_memory_mem_ck                      : out   std_logic_vector(0 downto 0);                     --                               .mem_ck
		ddr2_top_memory_mem_ck_n                    : out   std_logic_vector(0 downto 0);                     --                               .mem_ck_n
		ddr2_top_memory_mem_cke                     : out   std_logic_vector(0 downto 0);                     --                               .mem_cke
		ddr2_top_memory_mem_cs_n                    : out   std_logic_vector(0 downto 0);                     --                               .mem_cs_n
		ddr2_top_memory_mem_dm                      : out   std_logic_vector(3 downto 0);                     --                               .mem_dm
		ddr2_top_memory_mem_dq                      : inout std_logic_vector(31 downto 0) := (others => '0'); --                               .mem_dq
		ddr2_top_memory_mem_dqs                     : inout std_logic_vector(3 downto 0)  := (others => '0'); --                               .mem_dqs
		ddr2_top_memory_mem_dqs_n                   : inout std_logic_vector(3 downto 0)  := (others => '0'); --                               .mem_dqs_n
		ddr2_top_oct_rzqin                          : in    std_logic                     := '0';             --                   ddr2_top_oct.rzqin
		ddr2_top_status_local_init_done             : out   std_logic;                                        --                ddr2_top_status.local_init_done
		ddr2_top_status_local_cal_success           : out   std_logic;                                        --                               .local_cal_success
		ddr2_top_status_local_cal_fail              : out   std_logic;                                        --                               .local_cal_fail
		emac_gmii_connection_gmii_rx_d              : in    std_logic_vector(7 downto 0)  := (others => '0'); --           emac_gmii_connection.gmii_rx_d
		emac_gmii_connection_gmii_rx_dv             : in    std_logic                     := '0';             --                               .gmii_rx_dv
		emac_gmii_connection_gmii_rx_err            : in    std_logic                     := '0';             --                               .gmii_rx_err
		emac_gmii_connection_gmii_tx_d              : out   std_logic_vector(7 downto 0);                     --                               .gmii_tx_d
		emac_gmii_connection_gmii_tx_en             : out   std_logic;                                        --                               .gmii_tx_en
		emac_gmii_connection_gmii_tx_err            : out   std_logic;                                        --                               .gmii_tx_err
		emac_mdio_connection_mdc                    : out   std_logic;                                        --           emac_mdio_connection.mdc
		emac_mdio_connection_mdio_in                : in    std_logic                     := '0';             --                               .mdio_in
		emac_mdio_connection_mdio_out               : out   std_logic;                                        --                               .mdio_out
		emac_mdio_connection_mdio_oen               : out   std_logic;                                        --                               .mdio_oen
		emac_mii_connection_mii_rx_d                : in    std_logic_vector(3 downto 0)  := (others => '0'); --            emac_mii_connection.mii_rx_d
		emac_mii_connection_mii_rx_dv               : in    std_logic                     := '0';             --                               .mii_rx_dv
		emac_mii_connection_mii_rx_err              : in    std_logic                     := '0';             --                               .mii_rx_err
		emac_mii_connection_mii_tx_d                : out   std_logic_vector(3 downto 0);                     --                               .mii_tx_d
		emac_mii_connection_mii_tx_en               : out   std_logic;                                        --                               .mii_tx_en
		emac_mii_connection_mii_tx_err              : out   std_logic;                                        --                               .mii_tx_err
		emac_mii_connection_mii_crs                 : in    std_logic                     := '0';             --                               .mii_crs
		emac_mii_connection_mii_col                 : in    std_logic                     := '0';             --                               .mii_col
		emac_misc_connection_xon_gen                : in    std_logic                     := '0';             --           emac_misc_connection.xon_gen
		emac_misc_connection_xoff_gen               : in    std_logic                     := '0';             --                               .xoff_gen
		emac_misc_connection_ff_tx_crc_fwd          : in    std_logic                     := '0';             --                               .ff_tx_crc_fwd
		emac_misc_connection_ff_tx_septy            : out   std_logic;                                        --                               .ff_tx_septy
		emac_misc_connection_tx_ff_uflow            : out   std_logic;                                        --                               .tx_ff_uflow
		emac_misc_connection_ff_tx_a_full           : out   std_logic;                                        --                               .ff_tx_a_full
		emac_misc_connection_ff_tx_a_empty          : out   std_logic;                                        --                               .ff_tx_a_empty
		emac_misc_connection_rx_err_stat            : out   std_logic_vector(17 downto 0);                    --                               .rx_err_stat
		emac_misc_connection_rx_frm_type            : out   std_logic_vector(3 downto 0);                     --                               .rx_frm_type
		emac_misc_connection_ff_rx_dsav             : out   std_logic;                                        --                               .ff_rx_dsav
		emac_misc_connection_ff_rx_a_full           : out   std_logic;                                        --                               .ff_rx_a_full
		emac_misc_connection_ff_rx_a_empty          : out   std_logic;                                        --                               .ff_rx_a_empty
		emac_rx_clock_clk                           : in    std_logic                     := '0';             --                  emac_rx_clock.clk
		emac_status_connection_set_10               : in    std_logic                     := '0';             --         emac_status_connection.set_10
		emac_status_connection_set_1000             : in    std_logic                     := '0';             --                               .set_1000
		emac_status_connection_eth_mode             : out   std_logic;                                        --                               .eth_mode
		emac_status_connection_ena_10               : out   std_logic;                                        --                               .ena_10
		emac_tx_clock_clk                           : in    std_logic                     := '0';             --                  emac_tx_clock.clk
		enet_pll_clk125_clk                         : out   std_logic;                                        --                enet_pll_clk125.clk
		enet_pll_clk25_clk                          : out   std_logic;                                        --                 enet_pll_clk25.clk
		enet_pll_clk2_5_clk                         : out   std_logic;                                        --                enet_pll_clk2_5.clk
		enet_pll_locked_export                      : out   std_logic;                                        --                enet_pll_locked.export
		enet_pll_reset_reset                        : in    std_logic                     := '0';             --                 enet_pll_reset.reset
		led_pio_external_connection_export          : out   std_logic_vector(7 downto 0);                     --    led_pio_external_connection.export
		sdram_pll_sharing_pll_mem_clk               : out   std_logic;                                        --              sdram_pll_sharing.pll_mem_clk
		sdram_pll_sharing_pll_write_clk             : out   std_logic;                                        --                               .pll_write_clk
		sdram_pll_sharing_pll_locked                : out   std_logic;                                        --                               .pll_locked
		sdram_pll_sharing_pll_write_clk_pre_phy_clk : out   std_logic;                                        --                               .pll_write_clk_pre_phy_clk
		sdram_pll_sharing_pll_addr_cmd_clk          : out   std_logic;                                        --                               .pll_addr_cmd_clk
		sdram_pll_sharing_pll_avl_clk               : out   std_logic;                                        --                               .pll_avl_clk
		sdram_pll_sharing_pll_config_clk            : out   std_logic;                                        --                               .pll_config_clk
		sdram_pll_sharing_pll_mem_phy_clk           : out   std_logic;                                        --                               .pll_mem_phy_clk
		sdram_pll_sharing_afi_phy_clk               : out   std_logic;                                        --                               .afi_phy_clk
		sdram_pll_sharing_pll_avl_phy_clk           : out   std_logic                                         --                               .pll_avl_phy_clk
	);
end entity eth_std_main_system;

architecture rtl of eth_std_main_system is
	component eth_std_main_system_cpu is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(30 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(30 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component eth_std_main_system_cpu;

	component eth_std_main_system_enet_pll is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			outclk_1 : out std_logic;        -- clk
			outclk_2 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component eth_std_main_system_enet_pll;

	component eth_std_main_system_ethernet_subsystem is
		port (
			descriptor_memory_s2_address     : in  std_logic_vector(10 downto 0) := (others => 'X'); -- address
			descriptor_memory_s2_chipselect  : in  std_logic                     := 'X';             -- chipselect
			descriptor_memory_s2_clken       : in  std_logic                     := 'X';             -- clken
			descriptor_memory_s2_write       : in  std_logic                     := 'X';             -- write
			descriptor_memory_s2_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			descriptor_memory_s2_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			descriptor_memory_s2_byteenable  : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			ethernet_bridge_s0_waitrequest   : out std_logic;                                        -- waitrequest
			ethernet_bridge_s0_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			ethernet_bridge_s0_readdatavalid : out std_logic;                                        -- readdatavalid
			ethernet_bridge_s0_burstcount    : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			ethernet_bridge_s0_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			ethernet_bridge_s0_address       : in  std_logic_vector(10 downto 0) := (others => 'X'); -- address
			ethernet_bridge_s0_write         : in  std_logic                     := 'X';             -- write
			ethernet_bridge_s0_read          : in  std_logic                     := 'X';             -- read
			ethernet_bridge_s0_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			ethernet_bridge_s0_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			ethernet_subsys_clk_in_clk       : in  std_logic                     := 'X';             -- clk
			ethernet_subsys_reset_in_reset_n : in  std_logic                     := 'X';             -- reset_n
			mac_gmii_connection_gmii_rx_d    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- gmii_rx_d
			mac_gmii_connection_gmii_rx_dv   : in  std_logic                     := 'X';             -- gmii_rx_dv
			mac_gmii_connection_gmii_rx_err  : in  std_logic                     := 'X';             -- gmii_rx_err
			mac_gmii_connection_gmii_tx_d    : out std_logic_vector(7 downto 0);                     -- gmii_tx_d
			mac_gmii_connection_gmii_tx_en   : out std_logic;                                        -- gmii_tx_en
			mac_gmii_connection_gmii_tx_err  : out std_logic;                                        -- gmii_tx_err
			mac_mdio_connection_mdc          : out std_logic;                                        -- mdc
			mac_mdio_connection_mdio_in      : in  std_logic                     := 'X';             -- mdio_in
			mac_mdio_connection_mdio_out     : out std_logic;                                        -- mdio_out
			mac_mdio_connection_mdio_oen     : out std_logic;                                        -- mdio_oen
			mac_mii_connection_mii_rx_d      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- mii_rx_d
			mac_mii_connection_mii_rx_dv     : in  std_logic                     := 'X';             -- mii_rx_dv
			mac_mii_connection_mii_rx_err    : in  std_logic                     := 'X';             -- mii_rx_err
			mac_mii_connection_mii_tx_d      : out std_logic_vector(3 downto 0);                     -- mii_tx_d
			mac_mii_connection_mii_tx_en     : out std_logic;                                        -- mii_tx_en
			mac_mii_connection_mii_tx_err    : out std_logic;                                        -- mii_tx_err
			mac_mii_connection_mii_crs       : in  std_logic                     := 'X';             -- mii_crs
			mac_mii_connection_mii_col       : in  std_logic                     := 'X';             -- mii_col
			mac_status_connection_set_10     : in  std_logic                     := 'X';             -- set_10
			mac_status_connection_set_1000   : in  std_logic                     := 'X';             -- set_1000
			mac_status_connection_eth_mode   : out std_logic;                                        -- eth_mode
			mac_status_connection_ena_10     : out std_logic;                                        -- ena_10
			misc_connection_xon_gen          : in  std_logic                     := 'X';             -- xon_gen
			misc_connection_xoff_gen         : in  std_logic                     := 'X';             -- xoff_gen
			misc_connection_ff_tx_crc_fwd    : in  std_logic                     := 'X';             -- ff_tx_crc_fwd
			misc_connection_ff_tx_septy      : out std_logic;                                        -- ff_tx_septy
			misc_connection_tx_ff_uflow      : out std_logic;                                        -- tx_ff_uflow
			misc_connection_ff_tx_a_full     : out std_logic;                                        -- ff_tx_a_full
			misc_connection_ff_tx_a_empty    : out std_logic;                                        -- ff_tx_a_empty
			misc_connection_rx_err_stat      : out std_logic_vector(17 downto 0);                    -- rx_err_stat
			misc_connection_rx_frm_type      : out std_logic_vector(3 downto 0);                     -- rx_frm_type
			misc_connection_ff_rx_dsav       : out std_logic;                                        -- ff_rx_dsav
			misc_connection_ff_rx_a_full     : out std_logic;                                        -- ff_rx_a_full
			misc_connection_ff_rx_a_empty    : out std_logic;                                        -- ff_rx_a_empty
			rx_clock_clk                     : in  std_logic                     := 'X';             -- clk
			sgdma_bridge_m0_waitrequest      : in  std_logic                     := 'X';             -- waitrequest
			sgdma_bridge_m0_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sgdma_bridge_m0_readdatavalid    : in  std_logic                     := 'X';             -- readdatavalid
			sgdma_bridge_m0_burstcount       : out std_logic_vector(0 downto 0);                     -- burstcount
			sgdma_bridge_m0_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			sgdma_bridge_m0_address          : out std_logic_vector(30 downto 0);                    -- address
			sgdma_bridge_m0_write            : out std_logic;                                        -- write
			sgdma_bridge_m0_read             : out std_logic;                                        -- read
			sgdma_bridge_m0_byteenable       : out std_logic_vector(3 downto 0);                     -- byteenable
			sgdma_bridge_m0_debugaccess      : out std_logic;                                        -- debugaccess
			sgdma_rx_csr_irq_irq             : out std_logic;                                        -- irq
			sgdma_tx_csr_irq_irq             : out std_logic;                                        -- irq
			tx_clock_clk                     : in  std_logic                     := 'X'              -- clk
		);
	end component eth_std_main_system_ethernet_subsystem;

	component eth_std_main_system_peripheral_subsystem is
		port (
			button_pio_external_connection_export : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- export
			button_pio_irq_irq                    : out std_logic;                                        -- irq
			high_res_timer_irq_irq                : out std_logic;                                        -- irq
			jtag_uart_irq_irq                     : out std_logic;                                        -- irq
			led_pio_external_connection_export    : out std_logic_vector(7 downto 0);                     -- export
			peripheral_bridge_s0_waitrequest      : out std_logic;                                        -- waitrequest
			peripheral_bridge_s0_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			peripheral_bridge_s0_readdatavalid    : out std_logic;                                        -- readdatavalid
			peripheral_bridge_s0_burstcount       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			peripheral_bridge_s0_writedata        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			peripheral_bridge_s0_address          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			peripheral_bridge_s0_write            : in  std_logic                     := 'X';             -- write
			peripheral_bridge_s0_read             : in  std_logic                     := 'X';             -- read
			peripheral_bridge_s0_byteenable       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			peripheral_bridge_s0_debugaccess      : in  std_logic                     := 'X';             -- debugaccess
			peripheral_subsys_clk_in_clk          : in  std_logic                     := 'X';             -- clk
			peripheral_subsys_reset_in_reset_n    : in  std_logic                     := 'X';             -- reset_n
			sys_clk_timer_irq_irq                 : out std_logic                                         -- irq
		);
	end component eth_std_main_system_peripheral_subsystem;

	component eth_std_main_system_sdram is
		port (
			pll_ref_clk                : in    std_logic                     := 'X';             -- clk
			global_reset_n             : in    std_logic                     := 'X';             -- reset_n
			soft_reset_n               : in    std_logic                     := 'X';             -- reset_n
			afi_clk                    : out   std_logic;                                        -- clk
			afi_half_clk               : out   std_logic;                                        -- clk
			afi_reset_n                : out   std_logic;                                        -- reset_n
			afi_reset_export_n         : out   std_logic;                                        -- reset_n
			mem_ca                     : out   std_logic_vector(9 downto 0);                     -- mem_ca
			mem_ck                     : out   std_logic_vector(0 downto 0);                     -- mem_ck
			mem_ck_n                   : out   std_logic_vector(0 downto 0);                     -- mem_ck_n
			mem_cke                    : out   std_logic_vector(0 downto 0);                     -- mem_cke
			mem_cs_n                   : out   std_logic_vector(0 downto 0);                     -- mem_cs_n
			mem_dm                     : out   std_logic_vector(3 downto 0);                     -- mem_dm
			mem_dq                     : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs                    : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n                  : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			avl_ready_0                : out   std_logic;                                        -- waitrequest_n
			avl_burstbegin_0           : in    std_logic                     := 'X';             -- beginbursttransfer
			avl_addr_0                 : in    std_logic_vector(26 downto 0) := (others => 'X'); -- address
			avl_rdata_valid_0          : out   std_logic;                                        -- readdatavalid
			avl_rdata_0                : out   std_logic_vector(31 downto 0);                    -- readdata
			avl_wdata_0                : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avl_be_0                   : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avl_read_req_0             : in    std_logic                     := 'X';             -- read
			avl_write_req_0            : in    std_logic                     := 'X';             -- write
			avl_size_0                 : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			mp_cmd_clk_0_clk           : in    std_logic                     := 'X';             -- clk
			mp_cmd_reset_n_0_reset_n   : in    std_logic                     := 'X';             -- reset_n
			mp_rfifo_clk_0_clk         : in    std_logic                     := 'X';             -- clk
			mp_rfifo_reset_n_0_reset_n : in    std_logic                     := 'X';             -- reset_n
			mp_wfifo_clk_0_clk         : in    std_logic                     := 'X';             -- clk
			mp_wfifo_reset_n_0_reset_n : in    std_logic                     := 'X';             -- reset_n
			local_init_done            : out   std_logic;                                        -- local_init_done
			local_cal_success          : out   std_logic;                                        -- local_cal_success
			local_cal_fail             : out   std_logic;                                        -- local_cal_fail
			oct_rzqin                  : in    std_logic                     := 'X';             -- rzqin
			pll_mem_clk                : out   std_logic;                                        -- pll_mem_clk
			pll_write_clk              : out   std_logic;                                        -- pll_write_clk
			pll_locked                 : out   std_logic;                                        -- pll_locked
			pll_write_clk_pre_phy_clk  : out   std_logic;                                        -- pll_write_clk_pre_phy_clk
			pll_addr_cmd_clk           : out   std_logic;                                        -- pll_addr_cmd_clk
			pll_avl_clk                : out   std_logic;                                        -- pll_avl_clk
			pll_config_clk             : out   std_logic;                                        -- pll_config_clk
			pll_mem_phy_clk            : out   std_logic;                                        -- pll_mem_phy_clk
			afi_phy_clk                : out   std_logic;                                        -- afi_phy_clk
			pll_avl_phy_clk            : out   std_logic                                         -- pll_avl_phy_clk
		);
	end component eth_std_main_system_sdram;

	component eth_std_main_system_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component eth_std_main_system_sysid;

	component eth_std_main_system_mm_interconnect_0 is
		port (
			clk_125_clk_clk                                                         : in  std_logic                     := 'X';             -- clk
			clk_50_clk_clk                                                          : in  std_logic                     := 'X';             -- clk
			cpu_reset_reset_bridge_in_reset_reset                                   : in  std_logic                     := 'X';             -- reset
			ethernet_subsystem_ethernet_subsys_reset_in_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			sdram_avl_0_translator_reset_reset_bridge_in_reset_reset                : in  std_logic                     := 'X';             -- reset
			sdram_mp_cmd_reset_n_0_reset_bridge_in_reset_reset                      : in  std_logic                     := 'X';             -- reset
			sysid_reset_reset_bridge_in_reset_reset                                 : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                                                 : in  std_logic_vector(30 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest                                             : out std_logic;                                        -- waitrequest
			cpu_data_master_byteenable                                              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                                                    : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                                                : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_readdatavalid                                           : out std_logic;                                        -- readdatavalid
			cpu_data_master_write                                                   : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata                                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess                                             : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address                                          : in  std_logic_vector(30 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest                                      : out std_logic;                                        -- waitrequest
			cpu_instruction_master_read                                             : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata                                         : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_instruction_master_readdatavalid                                    : out std_logic;                                        -- readdatavalid
			ethernet_subsystem_sgdma_bridge_m0_address                              : in  std_logic_vector(30 downto 0) := (others => 'X'); -- address
			ethernet_subsystem_sgdma_bridge_m0_waitrequest                          : out std_logic;                                        -- waitrequest
			ethernet_subsystem_sgdma_bridge_m0_burstcount                           : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			ethernet_subsystem_sgdma_bridge_m0_byteenable                           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			ethernet_subsystem_sgdma_bridge_m0_read                                 : in  std_logic                     := 'X';             -- read
			ethernet_subsystem_sgdma_bridge_m0_readdata                             : out std_logic_vector(31 downto 0);                    -- readdata
			ethernet_subsystem_sgdma_bridge_m0_readdatavalid                        : out std_logic;                                        -- readdatavalid
			ethernet_subsystem_sgdma_bridge_m0_write                                : in  std_logic                     := 'X';             -- write
			ethernet_subsystem_sgdma_bridge_m0_writedata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			ethernet_subsystem_sgdma_bridge_m0_debugaccess                          : in  std_logic                     := 'X';             -- debugaccess
			cpu_debug_mem_slave_address                                             : out std_logic_vector(8 downto 0);                     -- address
			cpu_debug_mem_slave_write                                               : out std_logic;                                        -- write
			cpu_debug_mem_slave_read                                                : out std_logic;                                        -- read
			cpu_debug_mem_slave_readdata                                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_debug_mem_slave_writedata                                           : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_debug_mem_slave_byteenable                                          : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_debug_mem_slave_waitrequest                                         : in  std_logic                     := 'X';             -- waitrequest
			cpu_debug_mem_slave_debugaccess                                         : out std_logic;                                        -- debugaccess
			ethernet_subsystem_descriptor_memory_s2_address                         : out std_logic_vector(10 downto 0);                    -- address
			ethernet_subsystem_descriptor_memory_s2_write                           : out std_logic;                                        -- write
			ethernet_subsystem_descriptor_memory_s2_readdata                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ethernet_subsystem_descriptor_memory_s2_writedata                       : out std_logic_vector(31 downto 0);                    -- writedata
			ethernet_subsystem_descriptor_memory_s2_byteenable                      : out std_logic_vector(3 downto 0);                     -- byteenable
			ethernet_subsystem_descriptor_memory_s2_chipselect                      : out std_logic;                                        -- chipselect
			ethernet_subsystem_descriptor_memory_s2_clken                           : out std_logic;                                        -- clken
			ethernet_subsystem_ethernet_bridge_s0_address                           : out std_logic_vector(10 downto 0);                    -- address
			ethernet_subsystem_ethernet_bridge_s0_write                             : out std_logic;                                        -- write
			ethernet_subsystem_ethernet_bridge_s0_read                              : out std_logic;                                        -- read
			ethernet_subsystem_ethernet_bridge_s0_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ethernet_subsystem_ethernet_bridge_s0_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			ethernet_subsystem_ethernet_bridge_s0_burstcount                        : out std_logic_vector(0 downto 0);                     -- burstcount
			ethernet_subsystem_ethernet_bridge_s0_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			ethernet_subsystem_ethernet_bridge_s0_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			ethernet_subsystem_ethernet_bridge_s0_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			ethernet_subsystem_ethernet_bridge_s0_debugaccess                       : out std_logic;                                        -- debugaccess
			peripheral_subsystem_peripheral_bridge_s0_address                       : out std_logic_vector(7 downto 0);                     -- address
			peripheral_subsystem_peripheral_bridge_s0_write                         : out std_logic;                                        -- write
			peripheral_subsystem_peripheral_bridge_s0_read                          : out std_logic;                                        -- read
			peripheral_subsystem_peripheral_bridge_s0_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			peripheral_subsystem_peripheral_bridge_s0_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			peripheral_subsystem_peripheral_bridge_s0_burstcount                    : out std_logic_vector(0 downto 0);                     -- burstcount
			peripheral_subsystem_peripheral_bridge_s0_byteenable                    : out std_logic_vector(3 downto 0);                     -- byteenable
			peripheral_subsystem_peripheral_bridge_s0_readdatavalid                 : in  std_logic                     := 'X';             -- readdatavalid
			peripheral_subsystem_peripheral_bridge_s0_waitrequest                   : in  std_logic                     := 'X';             -- waitrequest
			peripheral_subsystem_peripheral_bridge_s0_debugaccess                   : out std_logic;                                        -- debugaccess
			sdram_avl_0_address                                                     : out std_logic_vector(26 downto 0);                    -- address
			sdram_avl_0_write                                                       : out std_logic;                                        -- write
			sdram_avl_0_read                                                        : out std_logic;                                        -- read
			sdram_avl_0_readdata                                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sdram_avl_0_writedata                                                   : out std_logic_vector(31 downto 0);                    -- writedata
			sdram_avl_0_beginbursttransfer                                          : out std_logic;                                        -- beginbursttransfer
			sdram_avl_0_burstcount                                                  : out std_logic_vector(2 downto 0);                     -- burstcount
			sdram_avl_0_byteenable                                                  : out std_logic_vector(3 downto 0);                     -- byteenable
			sdram_avl_0_readdatavalid                                               : in  std_logic                     := 'X';             -- readdatavalid
			sdram_avl_0_waitrequest                                                 : in  std_logic                     := 'X';             -- waitrequest
			sysid_control_slave_address                                             : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata                                            : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component eth_std_main_system_mm_interconnect_0;

	component eth_std_main_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			receiver5_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component eth_std_main_system_irq_mapper;

	component eth_std_main_system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_in2      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component eth_std_main_system_rst_controller;

	component eth_std_main_system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component eth_std_main_system_rst_controller_001;

	component eth_std_main_system_rst_controller_006 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component eth_std_main_system_rst_controller_006;

	signal cpu_data_master_readdata                                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_waitrequest                                               : std_logic;                     -- mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_debugaccess                                               : std_logic;                     -- cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	signal cpu_data_master_address                                                   : std_logic_vector(30 downto 0); -- cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	signal cpu_data_master_byteenable                                                : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	signal cpu_data_master_read                                                      : std_logic;                     -- cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	signal cpu_data_master_readdatavalid                                             : std_logic;                     -- mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	signal cpu_data_master_write                                                     : std_logic;                     -- cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	signal cpu_data_master_writedata                                                 : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	signal cpu_instruction_master_readdata                                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_waitrequest                                        : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                            : std_logic_vector(30 downto 0); -- cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	signal cpu_instruction_master_read                                               : std_logic;                     -- cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	signal cpu_instruction_master_readdatavalid                                      : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	signal ethernet_subsystem_sgdma_bridge_m0_waitrequest                            : std_logic;                     -- mm_interconnect_0:ethernet_subsystem_sgdma_bridge_m0_waitrequest -> ethernet_subsystem:sgdma_bridge_m0_waitrequest
	signal ethernet_subsystem_sgdma_bridge_m0_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:ethernet_subsystem_sgdma_bridge_m0_readdata -> ethernet_subsystem:sgdma_bridge_m0_readdata
	signal ethernet_subsystem_sgdma_bridge_m0_debugaccess                            : std_logic;                     -- ethernet_subsystem:sgdma_bridge_m0_debugaccess -> mm_interconnect_0:ethernet_subsystem_sgdma_bridge_m0_debugaccess
	signal ethernet_subsystem_sgdma_bridge_m0_address                                : std_logic_vector(30 downto 0); -- ethernet_subsystem:sgdma_bridge_m0_address -> mm_interconnect_0:ethernet_subsystem_sgdma_bridge_m0_address
	signal ethernet_subsystem_sgdma_bridge_m0_read                                   : std_logic;                     -- ethernet_subsystem:sgdma_bridge_m0_read -> mm_interconnect_0:ethernet_subsystem_sgdma_bridge_m0_read
	signal ethernet_subsystem_sgdma_bridge_m0_byteenable                             : std_logic_vector(3 downto 0);  -- ethernet_subsystem:sgdma_bridge_m0_byteenable -> mm_interconnect_0:ethernet_subsystem_sgdma_bridge_m0_byteenable
	signal ethernet_subsystem_sgdma_bridge_m0_readdatavalid                          : std_logic;                     -- mm_interconnect_0:ethernet_subsystem_sgdma_bridge_m0_readdatavalid -> ethernet_subsystem:sgdma_bridge_m0_readdatavalid
	signal ethernet_subsystem_sgdma_bridge_m0_writedata                              : std_logic_vector(31 downto 0); -- ethernet_subsystem:sgdma_bridge_m0_writedata -> mm_interconnect_0:ethernet_subsystem_sgdma_bridge_m0_writedata
	signal ethernet_subsystem_sgdma_bridge_m0_write                                  : std_logic;                     -- ethernet_subsystem:sgdma_bridge_m0_write -> mm_interconnect_0:ethernet_subsystem_sgdma_bridge_m0_write
	signal ethernet_subsystem_sgdma_bridge_m0_burstcount                             : std_logic_vector(0 downto 0);  -- ethernet_subsystem:sgdma_bridge_m0_burstcount -> mm_interconnect_0:ethernet_subsystem_sgdma_bridge_m0_burstcount
	signal mm_interconnect_0_sdram_avl_0_beginbursttransfer                          : std_logic;                     -- mm_interconnect_0:sdram_avl_0_beginbursttransfer -> sdram:avl_burstbegin_0
	signal mm_interconnect_0_sdram_avl_0_readdata                                    : std_logic_vector(31 downto 0); -- sdram:avl_rdata_0 -> mm_interconnect_0:sdram_avl_0_readdata
	signal sdram_avl_0_waitrequest                                                   : std_logic;                     -- sdram:avl_ready_0 -> sdram_avl_0_waitrequest:in
	signal mm_interconnect_0_sdram_avl_0_address                                     : std_logic_vector(26 downto 0); -- mm_interconnect_0:sdram_avl_0_address -> sdram:avl_addr_0
	signal mm_interconnect_0_sdram_avl_0_read                                        : std_logic;                     -- mm_interconnect_0:sdram_avl_0_read -> sdram:avl_read_req_0
	signal mm_interconnect_0_sdram_avl_0_byteenable                                  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:sdram_avl_0_byteenable -> sdram:avl_be_0
	signal mm_interconnect_0_sdram_avl_0_readdatavalid                               : std_logic;                     -- sdram:avl_rdata_valid_0 -> mm_interconnect_0:sdram_avl_0_readdatavalid
	signal mm_interconnect_0_sdram_avl_0_write                                       : std_logic;                     -- mm_interconnect_0:sdram_avl_0_write -> sdram:avl_write_req_0
	signal mm_interconnect_0_sdram_avl_0_writedata                                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:sdram_avl_0_writedata -> sdram:avl_wdata_0
	signal mm_interconnect_0_sdram_avl_0_burstcount                                  : std_logic_vector(2 downto 0);  -- mm_interconnect_0:sdram_avl_0_burstcount -> sdram:avl_size_0
	signal mm_interconnect_0_sysid_control_slave_readdata                            : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                             : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                            : std_logic_vector(31 downto 0); -- cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest                         : std_logic;                     -- cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess                         : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                             : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                                : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                               : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	signal mm_interconnect_0_ethernet_subsystem_descriptor_memory_s2_chipselect      : std_logic;                     -- mm_interconnect_0:ethernet_subsystem_descriptor_memory_s2_chipselect -> ethernet_subsystem:descriptor_memory_s2_chipselect
	signal mm_interconnect_0_ethernet_subsystem_descriptor_memory_s2_readdata        : std_logic_vector(31 downto 0); -- ethernet_subsystem:descriptor_memory_s2_readdata -> mm_interconnect_0:ethernet_subsystem_descriptor_memory_s2_readdata
	signal mm_interconnect_0_ethernet_subsystem_descriptor_memory_s2_address         : std_logic_vector(10 downto 0); -- mm_interconnect_0:ethernet_subsystem_descriptor_memory_s2_address -> ethernet_subsystem:descriptor_memory_s2_address
	signal mm_interconnect_0_ethernet_subsystem_descriptor_memory_s2_byteenable      : std_logic_vector(3 downto 0);  -- mm_interconnect_0:ethernet_subsystem_descriptor_memory_s2_byteenable -> ethernet_subsystem:descriptor_memory_s2_byteenable
	signal mm_interconnect_0_ethernet_subsystem_descriptor_memory_s2_write           : std_logic;                     -- mm_interconnect_0:ethernet_subsystem_descriptor_memory_s2_write -> ethernet_subsystem:descriptor_memory_s2_write
	signal mm_interconnect_0_ethernet_subsystem_descriptor_memory_s2_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:ethernet_subsystem_descriptor_memory_s2_writedata -> ethernet_subsystem:descriptor_memory_s2_writedata
	signal mm_interconnect_0_ethernet_subsystem_descriptor_memory_s2_clken           : std_logic;                     -- mm_interconnect_0:ethernet_subsystem_descriptor_memory_s2_clken -> ethernet_subsystem:descriptor_memory_s2_clken
	signal mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_readdata          : std_logic_vector(31 downto 0); -- ethernet_subsystem:ethernet_bridge_s0_readdata -> mm_interconnect_0:ethernet_subsystem_ethernet_bridge_s0_readdata
	signal mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_waitrequest       : std_logic;                     -- ethernet_subsystem:ethernet_bridge_s0_waitrequest -> mm_interconnect_0:ethernet_subsystem_ethernet_bridge_s0_waitrequest
	signal mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_debugaccess       : std_logic;                     -- mm_interconnect_0:ethernet_subsystem_ethernet_bridge_s0_debugaccess -> ethernet_subsystem:ethernet_bridge_s0_debugaccess
	signal mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_address           : std_logic_vector(10 downto 0); -- mm_interconnect_0:ethernet_subsystem_ethernet_bridge_s0_address -> ethernet_subsystem:ethernet_bridge_s0_address
	signal mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_read              : std_logic;                     -- mm_interconnect_0:ethernet_subsystem_ethernet_bridge_s0_read -> ethernet_subsystem:ethernet_bridge_s0_read
	signal mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_byteenable        : std_logic_vector(3 downto 0);  -- mm_interconnect_0:ethernet_subsystem_ethernet_bridge_s0_byteenable -> ethernet_subsystem:ethernet_bridge_s0_byteenable
	signal mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_readdatavalid     : std_logic;                     -- ethernet_subsystem:ethernet_bridge_s0_readdatavalid -> mm_interconnect_0:ethernet_subsystem_ethernet_bridge_s0_readdatavalid
	signal mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_write             : std_logic;                     -- mm_interconnect_0:ethernet_subsystem_ethernet_bridge_s0_write -> ethernet_subsystem:ethernet_bridge_s0_write
	signal mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:ethernet_subsystem_ethernet_bridge_s0_writedata -> ethernet_subsystem:ethernet_bridge_s0_writedata
	signal mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_burstcount        : std_logic_vector(0 downto 0);  -- mm_interconnect_0:ethernet_subsystem_ethernet_bridge_s0_burstcount -> ethernet_subsystem:ethernet_bridge_s0_burstcount
	signal mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_readdata      : std_logic_vector(31 downto 0); -- peripheral_subsystem:peripheral_bridge_s0_readdata -> mm_interconnect_0:peripheral_subsystem_peripheral_bridge_s0_readdata
	signal mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_waitrequest   : std_logic;                     -- peripheral_subsystem:peripheral_bridge_s0_waitrequest -> mm_interconnect_0:peripheral_subsystem_peripheral_bridge_s0_waitrequest
	signal mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_debugaccess   : std_logic;                     -- mm_interconnect_0:peripheral_subsystem_peripheral_bridge_s0_debugaccess -> peripheral_subsystem:peripheral_bridge_s0_debugaccess
	signal mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_address       : std_logic_vector(7 downto 0);  -- mm_interconnect_0:peripheral_subsystem_peripheral_bridge_s0_address -> peripheral_subsystem:peripheral_bridge_s0_address
	signal mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_read          : std_logic;                     -- mm_interconnect_0:peripheral_subsystem_peripheral_bridge_s0_read -> peripheral_subsystem:peripheral_bridge_s0_read
	signal mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_byteenable    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:peripheral_subsystem_peripheral_bridge_s0_byteenable -> peripheral_subsystem:peripheral_bridge_s0_byteenable
	signal mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_readdatavalid : std_logic;                     -- peripheral_subsystem:peripheral_bridge_s0_readdatavalid -> mm_interconnect_0:peripheral_subsystem_peripheral_bridge_s0_readdatavalid
	signal mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_write         : std_logic;                     -- mm_interconnect_0:peripheral_subsystem_peripheral_bridge_s0_write -> peripheral_subsystem:peripheral_bridge_s0_write
	signal mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:peripheral_subsystem_peripheral_bridge_s0_writedata -> peripheral_subsystem:peripheral_bridge_s0_writedata
	signal mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_burstcount    : std_logic_vector(0 downto 0);  -- mm_interconnect_0:peripheral_subsystem_peripheral_bridge_s0_burstcount -> peripheral_subsystem:peripheral_bridge_s0_burstcount
	signal irq_mapper_receiver0_irq                                                  : std_logic;                     -- peripheral_subsystem:button_pio_irq_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                  : std_logic;                     -- peripheral_subsystem:high_res_timer_irq_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                                  : std_logic;                     -- peripheral_subsystem:jtag_uart_irq_irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                                  : std_logic;                     -- ethernet_subsystem:sgdma_rx_csr_irq_irq -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                                  : std_logic;                     -- ethernet_subsystem:sgdma_tx_csr_irq_irq -> irq_mapper:receiver4_irq
	signal irq_mapper_receiver5_irq                                                  : std_logic;                     -- peripheral_subsystem:sys_clk_timer_irq_irq -> irq_mapper:receiver5_irq
	signal cpu_irq_irq                                                               : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:irq
	signal rst_controller_reset_out_reset                                            : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal rst_controller_reset_out_reset_req                                        : std_logic;                     -- rst_controller:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	signal cpu_debug_reset_request_reset                                             : std_logic;                     -- cpu:debug_reset_request -> rst_controller:reset_in2
	signal rst_controller_001_reset_out_reset                                        : std_logic;                     -- rst_controller_001:reset_out -> rst_controller_001_reset_out_reset:in
	signal rst_controller_002_reset_out_reset                                        : std_logic;                     -- rst_controller_002:reset_out -> rst_controller_002_reset_out_reset:in
	signal rst_controller_003_reset_out_reset                                        : std_logic;                     -- rst_controller_003:reset_out -> rst_controller_003_reset_out_reset:in
	signal rst_controller_004_reset_out_reset                                        : std_logic;                     -- rst_controller_004:reset_out -> rst_controller_004_reset_out_reset:in
	signal rst_controller_005_reset_out_reset                                        : std_logic;                     -- rst_controller_005:reset_out -> [mm_interconnect_0:ethernet_subsystem_ethernet_subsys_reset_in_reset_bridge_in_reset_reset, mm_interconnect_0:sysid_reset_reset_bridge_in_reset_reset, rst_controller_005_reset_out_reset:in]
	signal rst_controller_006_reset_out_reset                                        : std_logic;                     -- rst_controller_006:reset_out -> [mm_interconnect_0:sdram_avl_0_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:sdram_mp_cmd_reset_n_0_reset_bridge_in_reset_reset]
	signal clk_125_clk_in_reset_reset_n_ports_inv                                    : std_logic;                     -- clk_125_clk_in_reset_reset_n:inv -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in1, rst_controller_004:reset_in1, rst_controller_005:reset_in1, rst_controller_006:reset_in0]
	signal clk_50_clk_in_reset_reset_n_ports_inv                                     : std_logic;                     -- clk_50_clk_in_reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0, rst_controller_004:reset_in0, rst_controller_005:reset_in0]
	signal mm_interconnect_0_sdram_avl_0_inv                                         : std_logic;                     -- sdram_avl_0_waitrequest:inv -> mm_interconnect_0:sdram_avl_0_waitrequest
	signal rst_controller_reset_out_reset_ports_inv                                  : std_logic;                     -- rst_controller_reset_out_reset:inv -> cpu:reset_n
	signal rst_controller_001_reset_out_reset_ports_inv                              : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> ethernet_subsystem:ethernet_subsys_reset_in_reset_n
	signal rst_controller_002_reset_out_reset_ports_inv                              : std_logic;                     -- rst_controller_002_reset_out_reset:inv -> peripheral_subsystem:peripheral_subsys_reset_in_reset_n
	signal rst_controller_003_reset_out_reset_ports_inv                              : std_logic;                     -- rst_controller_003_reset_out_reset:inv -> sdram:global_reset_n
	signal rst_controller_004_reset_out_reset_ports_inv                              : std_logic;                     -- rst_controller_004_reset_out_reset:inv -> sdram:soft_reset_n
	signal rst_controller_005_reset_out_reset_ports_inv                              : std_logic;                     -- rst_controller_005_reset_out_reset:inv -> sysid:reset_n

begin

	cpu : component eth_std_main_system_cpu
		port map (
			clk                                 => clk_50_clk_in_clk,                                 --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,          --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			d_readdatavalid                     => cpu_data_master_readdatavalid,                     --                          .readdatavalid
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			i_readdatavalid                     => cpu_instruction_master_readdatavalid,              --                          .readdatavalid
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	enet_pll : component eth_std_main_system_enet_pll
		port map (
			refclk   => clk_50_clk_in_clk,      --  refclk.clk
			rst      => enet_pll_reset_reset,   --   reset.reset
			outclk_0 => enet_pll_clk125_clk,    -- outclk0.clk
			outclk_1 => enet_pll_clk25_clk,     -- outclk1.clk
			outclk_2 => enet_pll_clk2_5_clk,    -- outclk2.clk
			locked   => enet_pll_locked_export  --  locked.export
		);

	ethernet_subsystem : component eth_std_main_system_ethernet_subsystem
		port map (
			descriptor_memory_s2_address     => mm_interconnect_0_ethernet_subsystem_descriptor_memory_s2_address,     --     descriptor_memory_s2.address
			descriptor_memory_s2_chipselect  => mm_interconnect_0_ethernet_subsystem_descriptor_memory_s2_chipselect,  --                         .chipselect
			descriptor_memory_s2_clken       => mm_interconnect_0_ethernet_subsystem_descriptor_memory_s2_clken,       --                         .clken
			descriptor_memory_s2_write       => mm_interconnect_0_ethernet_subsystem_descriptor_memory_s2_write,       --                         .write
			descriptor_memory_s2_readdata    => mm_interconnect_0_ethernet_subsystem_descriptor_memory_s2_readdata,    --                         .readdata
			descriptor_memory_s2_writedata   => mm_interconnect_0_ethernet_subsystem_descriptor_memory_s2_writedata,   --                         .writedata
			descriptor_memory_s2_byteenable  => mm_interconnect_0_ethernet_subsystem_descriptor_memory_s2_byteenable,  --                         .byteenable
			ethernet_bridge_s0_waitrequest   => mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_waitrequest,   --       ethernet_bridge_s0.waitrequest
			ethernet_bridge_s0_readdata      => mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_readdata,      --                         .readdata
			ethernet_bridge_s0_readdatavalid => mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_readdatavalid, --                         .readdatavalid
			ethernet_bridge_s0_burstcount    => mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_burstcount,    --                         .burstcount
			ethernet_bridge_s0_writedata     => mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_writedata,     --                         .writedata
			ethernet_bridge_s0_address       => mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_address,       --                         .address
			ethernet_bridge_s0_write         => mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_write,         --                         .write
			ethernet_bridge_s0_read          => mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_read,          --                         .read
			ethernet_bridge_s0_byteenable    => mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_byteenable,    --                         .byteenable
			ethernet_bridge_s0_debugaccess   => mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_debugaccess,   --                         .debugaccess
			ethernet_subsys_clk_in_clk       => clk_50_clk_in_clk,                                                     --   ethernet_subsys_clk_in.clk
			ethernet_subsys_reset_in_reset_n => rst_controller_001_reset_out_reset_ports_inv,                          -- ethernet_subsys_reset_in.reset_n
			mac_gmii_connection_gmii_rx_d    => emac_gmii_connection_gmii_rx_d,                                        --      mac_gmii_connection.gmii_rx_d
			mac_gmii_connection_gmii_rx_dv   => emac_gmii_connection_gmii_rx_dv,                                       --                         .gmii_rx_dv
			mac_gmii_connection_gmii_rx_err  => emac_gmii_connection_gmii_rx_err,                                      --                         .gmii_rx_err
			mac_gmii_connection_gmii_tx_d    => emac_gmii_connection_gmii_tx_d,                                        --                         .gmii_tx_d
			mac_gmii_connection_gmii_tx_en   => emac_gmii_connection_gmii_tx_en,                                       --                         .gmii_tx_en
			mac_gmii_connection_gmii_tx_err  => emac_gmii_connection_gmii_tx_err,                                      --                         .gmii_tx_err
			mac_mdio_connection_mdc          => emac_mdio_connection_mdc,                                              --      mac_mdio_connection.mdc
			mac_mdio_connection_mdio_in      => emac_mdio_connection_mdio_in,                                          --                         .mdio_in
			mac_mdio_connection_mdio_out     => emac_mdio_connection_mdio_out,                                         --                         .mdio_out
			mac_mdio_connection_mdio_oen     => emac_mdio_connection_mdio_oen,                                         --                         .mdio_oen
			mac_mii_connection_mii_rx_d      => emac_mii_connection_mii_rx_d,                                          --       mac_mii_connection.mii_rx_d
			mac_mii_connection_mii_rx_dv     => emac_mii_connection_mii_rx_dv,                                         --                         .mii_rx_dv
			mac_mii_connection_mii_rx_err    => emac_mii_connection_mii_rx_err,                                        --                         .mii_rx_err
			mac_mii_connection_mii_tx_d      => emac_mii_connection_mii_tx_d,                                          --                         .mii_tx_d
			mac_mii_connection_mii_tx_en     => emac_mii_connection_mii_tx_en,                                         --                         .mii_tx_en
			mac_mii_connection_mii_tx_err    => emac_mii_connection_mii_tx_err,                                        --                         .mii_tx_err
			mac_mii_connection_mii_crs       => emac_mii_connection_mii_crs,                                           --                         .mii_crs
			mac_mii_connection_mii_col       => emac_mii_connection_mii_col,                                           --                         .mii_col
			mac_status_connection_set_10     => emac_status_connection_set_10,                                         --    mac_status_connection.set_10
			mac_status_connection_set_1000   => emac_status_connection_set_1000,                                       --                         .set_1000
			mac_status_connection_eth_mode   => emac_status_connection_eth_mode,                                       --                         .eth_mode
			mac_status_connection_ena_10     => emac_status_connection_ena_10,                                         --                         .ena_10
			misc_connection_xon_gen          => emac_misc_connection_xon_gen,                                          --          misc_connection.xon_gen
			misc_connection_xoff_gen         => emac_misc_connection_xoff_gen,                                         --                         .xoff_gen
			misc_connection_ff_tx_crc_fwd    => emac_misc_connection_ff_tx_crc_fwd,                                    --                         .ff_tx_crc_fwd
			misc_connection_ff_tx_septy      => emac_misc_connection_ff_tx_septy,                                      --                         .ff_tx_septy
			misc_connection_tx_ff_uflow      => emac_misc_connection_tx_ff_uflow,                                      --                         .tx_ff_uflow
			misc_connection_ff_tx_a_full     => emac_misc_connection_ff_tx_a_full,                                     --                         .ff_tx_a_full
			misc_connection_ff_tx_a_empty    => emac_misc_connection_ff_tx_a_empty,                                    --                         .ff_tx_a_empty
			misc_connection_rx_err_stat      => emac_misc_connection_rx_err_stat,                                      --                         .rx_err_stat
			misc_connection_rx_frm_type      => emac_misc_connection_rx_frm_type,                                      --                         .rx_frm_type
			misc_connection_ff_rx_dsav       => emac_misc_connection_ff_rx_dsav,                                       --                         .ff_rx_dsav
			misc_connection_ff_rx_a_full     => emac_misc_connection_ff_rx_a_full,                                     --                         .ff_rx_a_full
			misc_connection_ff_rx_a_empty    => emac_misc_connection_ff_rx_a_empty,                                    --                         .ff_rx_a_empty
			rx_clock_clk                     => emac_rx_clock_clk,                                                     --                 rx_clock.clk
			sgdma_bridge_m0_waitrequest      => ethernet_subsystem_sgdma_bridge_m0_waitrequest,                        --          sgdma_bridge_m0.waitrequest
			sgdma_bridge_m0_readdata         => ethernet_subsystem_sgdma_bridge_m0_readdata,                           --                         .readdata
			sgdma_bridge_m0_readdatavalid    => ethernet_subsystem_sgdma_bridge_m0_readdatavalid,                      --                         .readdatavalid
			sgdma_bridge_m0_burstcount       => ethernet_subsystem_sgdma_bridge_m0_burstcount,                         --                         .burstcount
			sgdma_bridge_m0_writedata        => ethernet_subsystem_sgdma_bridge_m0_writedata,                          --                         .writedata
			sgdma_bridge_m0_address          => ethernet_subsystem_sgdma_bridge_m0_address,                            --                         .address
			sgdma_bridge_m0_write            => ethernet_subsystem_sgdma_bridge_m0_write,                              --                         .write
			sgdma_bridge_m0_read             => ethernet_subsystem_sgdma_bridge_m0_read,                               --                         .read
			sgdma_bridge_m0_byteenable       => ethernet_subsystem_sgdma_bridge_m0_byteenable,                         --                         .byteenable
			sgdma_bridge_m0_debugaccess      => ethernet_subsystem_sgdma_bridge_m0_debugaccess,                        --                         .debugaccess
			sgdma_rx_csr_irq_irq             => irq_mapper_receiver3_irq,                                              --         sgdma_rx_csr_irq.irq
			sgdma_tx_csr_irq_irq             => irq_mapper_receiver4_irq,                                              --         sgdma_tx_csr_irq.irq
			tx_clock_clk                     => emac_tx_clock_clk                                                      --                 tx_clock.clk
		);

	peripheral_subsystem : component eth_std_main_system_peripheral_subsystem
		port map (
			button_pio_external_connection_export => button_pio_external_connection_export,                                     -- button_pio_external_connection.export
			button_pio_irq_irq                    => irq_mapper_receiver0_irq,                                                  --                 button_pio_irq.irq
			high_res_timer_irq_irq                => irq_mapper_receiver1_irq,                                                  --             high_res_timer_irq.irq
			jtag_uart_irq_irq                     => irq_mapper_receiver2_irq,                                                  --                  jtag_uart_irq.irq
			led_pio_external_connection_export    => led_pio_external_connection_export,                                        --    led_pio_external_connection.export
			peripheral_bridge_s0_waitrequest      => mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_waitrequest,   --           peripheral_bridge_s0.waitrequest
			peripheral_bridge_s0_readdata         => mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_readdata,      --                               .readdata
			peripheral_bridge_s0_readdatavalid    => mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_readdatavalid, --                               .readdatavalid
			peripheral_bridge_s0_burstcount       => mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_burstcount,    --                               .burstcount
			peripheral_bridge_s0_writedata        => mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_writedata,     --                               .writedata
			peripheral_bridge_s0_address          => mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_address,       --                               .address
			peripheral_bridge_s0_write            => mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_write,         --                               .write
			peripheral_bridge_s0_read             => mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_read,          --                               .read
			peripheral_bridge_s0_byteenable       => mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_byteenable,    --                               .byteenable
			peripheral_bridge_s0_debugaccess      => mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_debugaccess,   --                               .debugaccess
			peripheral_subsys_clk_in_clk          => clk_50_clk_in_clk,                                                         --       peripheral_subsys_clk_in.clk
			peripheral_subsys_reset_in_reset_n    => rst_controller_002_reset_out_reset_ports_inv,                              --     peripheral_subsys_reset_in.reset_n
			sys_clk_timer_irq_irq                 => irq_mapper_receiver5_irq                                                   --              sys_clk_timer_irq.irq
		);

	sdram : component eth_std_main_system_sdram
		port map (
			pll_ref_clk                => clk_125_clk_in_clk,                               --        pll_ref_clk.clk
			global_reset_n             => rst_controller_003_reset_out_reset_ports_inv,     --       global_reset.reset_n
			soft_reset_n               => rst_controller_004_reset_out_reset_ports_inv,     --         soft_reset.reset_n
			afi_clk                    => open,                                             --            afi_clk.clk
			afi_half_clk               => open,                                             --       afi_half_clk.clk
			afi_reset_n                => open,                                             --          afi_reset.reset_n
			afi_reset_export_n         => open,                                             --   afi_reset_export.reset_n
			mem_ca                     => ddr2_top_memory_mem_ca,                           --             memory.mem_ca
			mem_ck                     => ddr2_top_memory_mem_ck,                           --                   .mem_ck
			mem_ck_n                   => ddr2_top_memory_mem_ck_n,                         --                   .mem_ck_n
			mem_cke                    => ddr2_top_memory_mem_cke,                          --                   .mem_cke
			mem_cs_n                   => ddr2_top_memory_mem_cs_n,                         --                   .mem_cs_n
			mem_dm                     => ddr2_top_memory_mem_dm,                           --                   .mem_dm
			mem_dq                     => ddr2_top_memory_mem_dq,                           --                   .mem_dq
			mem_dqs                    => ddr2_top_memory_mem_dqs,                          --                   .mem_dqs
			mem_dqs_n                  => ddr2_top_memory_mem_dqs_n,                        --                   .mem_dqs_n
			avl_ready_0                => sdram_avl_0_waitrequest,                          --              avl_0.waitrequest_n
			avl_burstbegin_0           => mm_interconnect_0_sdram_avl_0_beginbursttransfer, --                   .beginbursttransfer
			avl_addr_0                 => mm_interconnect_0_sdram_avl_0_address,            --                   .address
			avl_rdata_valid_0          => mm_interconnect_0_sdram_avl_0_readdatavalid,      --                   .readdatavalid
			avl_rdata_0                => mm_interconnect_0_sdram_avl_0_readdata,           --                   .readdata
			avl_wdata_0                => mm_interconnect_0_sdram_avl_0_writedata,          --                   .writedata
			avl_be_0                   => mm_interconnect_0_sdram_avl_0_byteenable,         --                   .byteenable
			avl_read_req_0             => mm_interconnect_0_sdram_avl_0_read,               --                   .read
			avl_write_req_0            => mm_interconnect_0_sdram_avl_0_write,              --                   .write
			avl_size_0                 => mm_interconnect_0_sdram_avl_0_burstcount,         --                   .burstcount
			mp_cmd_clk_0_clk           => clk_125_clk_in_clk,                               --       mp_cmd_clk_0.clk
			mp_cmd_reset_n_0_reset_n   => clk_125_clk_in_reset_reset_n,                     --   mp_cmd_reset_n_0.reset_n
			mp_rfifo_clk_0_clk         => clk_125_clk_in_clk,                               --     mp_rfifo_clk_0.clk
			mp_rfifo_reset_n_0_reset_n => clk_125_clk_in_reset_reset_n,                     -- mp_rfifo_reset_n_0.reset_n
			mp_wfifo_clk_0_clk         => clk_125_clk_in_clk,                               --     mp_wfifo_clk_0.clk
			mp_wfifo_reset_n_0_reset_n => clk_125_clk_in_reset_reset_n,                     -- mp_wfifo_reset_n_0.reset_n
			local_init_done            => ddr2_top_status_local_init_done,                  --             status.local_init_done
			local_cal_success          => ddr2_top_status_local_cal_success,                --                   .local_cal_success
			local_cal_fail             => ddr2_top_status_local_cal_fail,                   --                   .local_cal_fail
			oct_rzqin                  => ddr2_top_oct_rzqin,                               --                oct.rzqin
			pll_mem_clk                => sdram_pll_sharing_pll_mem_clk,                    --        pll_sharing.pll_mem_clk
			pll_write_clk              => sdram_pll_sharing_pll_write_clk,                  --                   .pll_write_clk
			pll_locked                 => sdram_pll_sharing_pll_locked,                     --                   .pll_locked
			pll_write_clk_pre_phy_clk  => sdram_pll_sharing_pll_write_clk_pre_phy_clk,      --                   .pll_write_clk_pre_phy_clk
			pll_addr_cmd_clk           => sdram_pll_sharing_pll_addr_cmd_clk,               --                   .pll_addr_cmd_clk
			pll_avl_clk                => sdram_pll_sharing_pll_avl_clk,                    --                   .pll_avl_clk
			pll_config_clk             => sdram_pll_sharing_pll_config_clk,                 --                   .pll_config_clk
			pll_mem_phy_clk            => sdram_pll_sharing_pll_mem_phy_clk,                --                   .pll_mem_phy_clk
			afi_phy_clk                => sdram_pll_sharing_afi_phy_clk,                    --                   .afi_phy_clk
			pll_avl_phy_clk            => sdram_pll_sharing_pll_avl_phy_clk                 --                   .pll_avl_phy_clk
		);

	sysid : component eth_std_main_system_sysid
		port map (
			clock    => clk_50_clk_in_clk,                                --           clk.clk
			reset_n  => rst_controller_005_reset_out_reset_ports_inv,     --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component eth_std_main_system_mm_interconnect_0
		port map (
			clk_125_clk_clk                                                         => clk_125_clk_in_clk,                                                        --                                                       clk_125_clk.clk
			clk_50_clk_clk                                                          => clk_50_clk_in_clk,                                                         --                                                        clk_50_clk.clk
			cpu_reset_reset_bridge_in_reset_reset                                   => rst_controller_reset_out_reset,                                            --                                   cpu_reset_reset_bridge_in_reset.reset
			ethernet_subsystem_ethernet_subsys_reset_in_reset_bridge_in_reset_reset => rst_controller_005_reset_out_reset,                                        -- ethernet_subsystem_ethernet_subsys_reset_in_reset_bridge_in_reset.reset
			sdram_avl_0_translator_reset_reset_bridge_in_reset_reset                => rst_controller_006_reset_out_reset,                                        --                sdram_avl_0_translator_reset_reset_bridge_in_reset.reset
			sdram_mp_cmd_reset_n_0_reset_bridge_in_reset_reset                      => rst_controller_006_reset_out_reset,                                        --                      sdram_mp_cmd_reset_n_0_reset_bridge_in_reset.reset
			sysid_reset_reset_bridge_in_reset_reset                                 => rst_controller_005_reset_out_reset,                                        --                                 sysid_reset_reset_bridge_in_reset.reset
			cpu_data_master_address                                                 => cpu_data_master_address,                                                   --                                                   cpu_data_master.address
			cpu_data_master_waitrequest                                             => cpu_data_master_waitrequest,                                               --                                                                  .waitrequest
			cpu_data_master_byteenable                                              => cpu_data_master_byteenable,                                                --                                                                  .byteenable
			cpu_data_master_read                                                    => cpu_data_master_read,                                                      --                                                                  .read
			cpu_data_master_readdata                                                => cpu_data_master_readdata,                                                  --                                                                  .readdata
			cpu_data_master_readdatavalid                                           => cpu_data_master_readdatavalid,                                             --                                                                  .readdatavalid
			cpu_data_master_write                                                   => cpu_data_master_write,                                                     --                                                                  .write
			cpu_data_master_writedata                                               => cpu_data_master_writedata,                                                 --                                                                  .writedata
			cpu_data_master_debugaccess                                             => cpu_data_master_debugaccess,                                               --                                                                  .debugaccess
			cpu_instruction_master_address                                          => cpu_instruction_master_address,                                            --                                            cpu_instruction_master.address
			cpu_instruction_master_waitrequest                                      => cpu_instruction_master_waitrequest,                                        --                                                                  .waitrequest
			cpu_instruction_master_read                                             => cpu_instruction_master_read,                                               --                                                                  .read
			cpu_instruction_master_readdata                                         => cpu_instruction_master_readdata,                                           --                                                                  .readdata
			cpu_instruction_master_readdatavalid                                    => cpu_instruction_master_readdatavalid,                                      --                                                                  .readdatavalid
			ethernet_subsystem_sgdma_bridge_m0_address                              => ethernet_subsystem_sgdma_bridge_m0_address,                                --                                ethernet_subsystem_sgdma_bridge_m0.address
			ethernet_subsystem_sgdma_bridge_m0_waitrequest                          => ethernet_subsystem_sgdma_bridge_m0_waitrequest,                            --                                                                  .waitrequest
			ethernet_subsystem_sgdma_bridge_m0_burstcount                           => ethernet_subsystem_sgdma_bridge_m0_burstcount,                             --                                                                  .burstcount
			ethernet_subsystem_sgdma_bridge_m0_byteenable                           => ethernet_subsystem_sgdma_bridge_m0_byteenable,                             --                                                                  .byteenable
			ethernet_subsystem_sgdma_bridge_m0_read                                 => ethernet_subsystem_sgdma_bridge_m0_read,                                   --                                                                  .read
			ethernet_subsystem_sgdma_bridge_m0_readdata                             => ethernet_subsystem_sgdma_bridge_m0_readdata,                               --                                                                  .readdata
			ethernet_subsystem_sgdma_bridge_m0_readdatavalid                        => ethernet_subsystem_sgdma_bridge_m0_readdatavalid,                          --                                                                  .readdatavalid
			ethernet_subsystem_sgdma_bridge_m0_write                                => ethernet_subsystem_sgdma_bridge_m0_write,                                  --                                                                  .write
			ethernet_subsystem_sgdma_bridge_m0_writedata                            => ethernet_subsystem_sgdma_bridge_m0_writedata,                              --                                                                  .writedata
			ethernet_subsystem_sgdma_bridge_m0_debugaccess                          => ethernet_subsystem_sgdma_bridge_m0_debugaccess,                            --                                                                  .debugaccess
			cpu_debug_mem_slave_address                                             => mm_interconnect_0_cpu_debug_mem_slave_address,                             --                                               cpu_debug_mem_slave.address
			cpu_debug_mem_slave_write                                               => mm_interconnect_0_cpu_debug_mem_slave_write,                               --                                                                  .write
			cpu_debug_mem_slave_read                                                => mm_interconnect_0_cpu_debug_mem_slave_read,                                --                                                                  .read
			cpu_debug_mem_slave_readdata                                            => mm_interconnect_0_cpu_debug_mem_slave_readdata,                            --                                                                  .readdata
			cpu_debug_mem_slave_writedata                                           => mm_interconnect_0_cpu_debug_mem_slave_writedata,                           --                                                                  .writedata
			cpu_debug_mem_slave_byteenable                                          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,                          --                                                                  .byteenable
			cpu_debug_mem_slave_waitrequest                                         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,                         --                                                                  .waitrequest
			cpu_debug_mem_slave_debugaccess                                         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,                         --                                                                  .debugaccess
			ethernet_subsystem_descriptor_memory_s2_address                         => mm_interconnect_0_ethernet_subsystem_descriptor_memory_s2_address,         --                           ethernet_subsystem_descriptor_memory_s2.address
			ethernet_subsystem_descriptor_memory_s2_write                           => mm_interconnect_0_ethernet_subsystem_descriptor_memory_s2_write,           --                                                                  .write
			ethernet_subsystem_descriptor_memory_s2_readdata                        => mm_interconnect_0_ethernet_subsystem_descriptor_memory_s2_readdata,        --                                                                  .readdata
			ethernet_subsystem_descriptor_memory_s2_writedata                       => mm_interconnect_0_ethernet_subsystem_descriptor_memory_s2_writedata,       --                                                                  .writedata
			ethernet_subsystem_descriptor_memory_s2_byteenable                      => mm_interconnect_0_ethernet_subsystem_descriptor_memory_s2_byteenable,      --                                                                  .byteenable
			ethernet_subsystem_descriptor_memory_s2_chipselect                      => mm_interconnect_0_ethernet_subsystem_descriptor_memory_s2_chipselect,      --                                                                  .chipselect
			ethernet_subsystem_descriptor_memory_s2_clken                           => mm_interconnect_0_ethernet_subsystem_descriptor_memory_s2_clken,           --                                                                  .clken
			ethernet_subsystem_ethernet_bridge_s0_address                           => mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_address,           --                             ethernet_subsystem_ethernet_bridge_s0.address
			ethernet_subsystem_ethernet_bridge_s0_write                             => mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_write,             --                                                                  .write
			ethernet_subsystem_ethernet_bridge_s0_read                              => mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_read,              --                                                                  .read
			ethernet_subsystem_ethernet_bridge_s0_readdata                          => mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_readdata,          --                                                                  .readdata
			ethernet_subsystem_ethernet_bridge_s0_writedata                         => mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_writedata,         --                                                                  .writedata
			ethernet_subsystem_ethernet_bridge_s0_burstcount                        => mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_burstcount,        --                                                                  .burstcount
			ethernet_subsystem_ethernet_bridge_s0_byteenable                        => mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_byteenable,        --                                                                  .byteenable
			ethernet_subsystem_ethernet_bridge_s0_readdatavalid                     => mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_readdatavalid,     --                                                                  .readdatavalid
			ethernet_subsystem_ethernet_bridge_s0_waitrequest                       => mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_waitrequest,       --                                                                  .waitrequest
			ethernet_subsystem_ethernet_bridge_s0_debugaccess                       => mm_interconnect_0_ethernet_subsystem_ethernet_bridge_s0_debugaccess,       --                                                                  .debugaccess
			peripheral_subsystem_peripheral_bridge_s0_address                       => mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_address,       --                         peripheral_subsystem_peripheral_bridge_s0.address
			peripheral_subsystem_peripheral_bridge_s0_write                         => mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_write,         --                                                                  .write
			peripheral_subsystem_peripheral_bridge_s0_read                          => mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_read,          --                                                                  .read
			peripheral_subsystem_peripheral_bridge_s0_readdata                      => mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_readdata,      --                                                                  .readdata
			peripheral_subsystem_peripheral_bridge_s0_writedata                     => mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_writedata,     --                                                                  .writedata
			peripheral_subsystem_peripheral_bridge_s0_burstcount                    => mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_burstcount,    --                                                                  .burstcount
			peripheral_subsystem_peripheral_bridge_s0_byteenable                    => mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_byteenable,    --                                                                  .byteenable
			peripheral_subsystem_peripheral_bridge_s0_readdatavalid                 => mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_readdatavalid, --                                                                  .readdatavalid
			peripheral_subsystem_peripheral_bridge_s0_waitrequest                   => mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_waitrequest,   --                                                                  .waitrequest
			peripheral_subsystem_peripheral_bridge_s0_debugaccess                   => mm_interconnect_0_peripheral_subsystem_peripheral_bridge_s0_debugaccess,   --                                                                  .debugaccess
			sdram_avl_0_address                                                     => mm_interconnect_0_sdram_avl_0_address,                                     --                                                       sdram_avl_0.address
			sdram_avl_0_write                                                       => mm_interconnect_0_sdram_avl_0_write,                                       --                                                                  .write
			sdram_avl_0_read                                                        => mm_interconnect_0_sdram_avl_0_read,                                        --                                                                  .read
			sdram_avl_0_readdata                                                    => mm_interconnect_0_sdram_avl_0_readdata,                                    --                                                                  .readdata
			sdram_avl_0_writedata                                                   => mm_interconnect_0_sdram_avl_0_writedata,                                   --                                                                  .writedata
			sdram_avl_0_beginbursttransfer                                          => mm_interconnect_0_sdram_avl_0_beginbursttransfer,                          --                                                                  .beginbursttransfer
			sdram_avl_0_burstcount                                                  => mm_interconnect_0_sdram_avl_0_burstcount,                                  --                                                                  .burstcount
			sdram_avl_0_byteenable                                                  => mm_interconnect_0_sdram_avl_0_byteenable,                                  --                                                                  .byteenable
			sdram_avl_0_readdatavalid                                               => mm_interconnect_0_sdram_avl_0_readdatavalid,                               --                                                                  .readdatavalid
			sdram_avl_0_waitrequest                                                 => mm_interconnect_0_sdram_avl_0_inv,                                         --                                                                  .waitrequest
			sysid_control_slave_address                                             => mm_interconnect_0_sysid_control_slave_address,                             --                                               sysid_control_slave.address
			sysid_control_slave_readdata                                            => mm_interconnect_0_sysid_control_slave_readdata                             --                                                                  .readdata
		);

	irq_mapper : component eth_std_main_system_irq_mapper
		port map (
			clk           => clk_50_clk_in_clk,              --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,       -- receiver4.irq
			receiver5_irq => irq_mapper_receiver5_irq,       -- receiver5.irq
			sender_irq    => cpu_irq_irq                     --    sender.irq
		);

	rst_controller : component eth_std_main_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 3,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => clk_50_clk_in_reset_reset_n_ports_inv,  -- reset_in0.reset
			reset_in1      => clk_125_clk_in_reset_reset_n_ports_inv, -- reset_in1.reset
			reset_in2      => cpu_debug_reset_request_reset,          -- reset_in2.reset
			clk            => clk_50_clk_in_clk,                      --       clk.clk
			reset_out      => rst_controller_reset_out_reset,         -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,     --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_001 : component eth_std_main_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => clk_50_clk_in_reset_reset_n_ports_inv,  -- reset_in0.reset
			reset_in1      => clk_125_clk_in_reset_reset_n_ports_inv, -- reset_in1.reset
			clk            => open,                                   --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => open,                                   -- (terminated)
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_002 : component eth_std_main_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => clk_50_clk_in_reset_reset_n_ports_inv,  -- reset_in0.reset
			reset_in1      => clk_125_clk_in_reset_reset_n_ports_inv, -- reset_in1.reset
			clk            => open,                                   --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,     -- reset_out.reset
			reset_req      => open,                                   -- (terminated)
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_003 : component eth_std_main_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => clk_50_clk_in_reset_reset_n_ports_inv,  -- reset_in0.reset
			reset_in1      => clk_125_clk_in_reset_reset_n_ports_inv, -- reset_in1.reset
			clk            => open,                                   --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset,     -- reset_out.reset
			reset_req      => open,                                   -- (terminated)
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_004 : component eth_std_main_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => clk_50_clk_in_reset_reset_n_ports_inv,  -- reset_in0.reset
			reset_in1      => clk_125_clk_in_reset_reset_n_ports_inv, -- reset_in1.reset
			clk            => open,                                   --       clk.clk
			reset_out      => rst_controller_004_reset_out_reset,     -- reset_out.reset
			reset_req      => open,                                   -- (terminated)
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_005 : component eth_std_main_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => clk_50_clk_in_reset_reset_n_ports_inv,  -- reset_in0.reset
			reset_in1      => clk_125_clk_in_reset_reset_n_ports_inv, -- reset_in1.reset
			clk            => clk_50_clk_in_clk,                      --       clk.clk
			reset_out      => rst_controller_005_reset_out_reset,     -- reset_out.reset
			reset_req      => open,                                   -- (terminated)
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_006 : component eth_std_main_system_rst_controller_006
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => clk_125_clk_in_reset_reset_n_ports_inv, -- reset_in0.reset
			clk            => clk_125_clk_in_clk,                     --       clk.clk
			reset_out      => rst_controller_006_reset_out_reset,     -- reset_out.reset
			reset_req      => open,                                   -- (terminated)
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	clk_125_clk_in_reset_reset_n_ports_inv <= not clk_125_clk_in_reset_reset_n;

	clk_50_clk_in_reset_reset_n_ports_inv <= not clk_50_clk_in_reset_reset_n;

	mm_interconnect_0_sdram_avl_0_inv <= not sdram_avl_0_waitrequest;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

	rst_controller_003_reset_out_reset_ports_inv <= not rst_controller_003_reset_out_reset;

	rst_controller_004_reset_out_reset_ports_inv <= not rst_controller_004_reset_out_reset;

	rst_controller_005_reset_out_reset_ports_inv <= not rst_controller_005_reset_out_reset;

end architecture rtl; -- of eth_std_main_system
